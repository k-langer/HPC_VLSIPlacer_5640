module mips ( gnd, vdd, clk, reset, instr, readdata, pc, memwrite, aluout, writedata);

input gnd, vdd;
input clk;
input reset;
output memwrite;
input [31:0] instr;
input [31:0] readdata;
output [31:0] pc;
output [31:0] aluout;
output [31:0] writedata;

	BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(pc_0__RAW), .Y(pc[0]) );
	BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(pc_1__RAW), .Y(pc[1]) );
	BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(pc_2__RAW), .Y(pc[2]) );
	BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(pc_3__RAW), .Y(pc[3]) );
	BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(pc_4__RAW), .Y(pc[4]) );
	BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(pc_5__RAW), .Y(pc[5]) );
	BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(pc_6__RAW), .Y(pc[6]) );
	BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(pc_7__RAW), .Y(pc[7]) );
	BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(pc_8__RAW), .Y(pc[8]) );
	BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(pc_9__RAW), .Y(pc[9]) );
	BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(pc_10__RAW), .Y(pc[10]) );
	BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(pc_11__RAW), .Y(pc[11]) );
	BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(pc_12__RAW), .Y(pc[12]) );
	BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(pc_13__RAW), .Y(pc[13]) );
	BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(pc_14__RAW), .Y(pc[14]) );
	BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(pc_15__RAW), .Y(pc[15]) );
	BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(pc_16__RAW), .Y(pc[16]) );
	BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(pc_17__RAW), .Y(pc[17]) );
	BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(pc_18__RAW), .Y(pc[18]) );
	BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(pc_19__RAW), .Y(pc[19]) );
	BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(pc_20__RAW), .Y(pc[20]) );
	BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(pc_21__RAW), .Y(pc[21]) );
	BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(pc_22__RAW), .Y(pc[22]) );
	BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(pc_23__RAW), .Y(pc[23]) );
	BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(pc_24__RAW), .Y(pc[24]) );
	BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(pc_25__RAW), .Y(pc[25]) );
	BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(pc_26__RAW), .Y(pc[26]) );
	BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(pc_27__RAW), .Y(pc[27]) );
	BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(pc_28__RAW), .Y(pc[28]) );
	BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(pc_29__RAW), .Y(pc[29]) );
	BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(pc_30__RAW), .Y(pc[30]) );
	BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(pc_31__RAW), .Y(pc[31]) );
	BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(memwrite_RAW), .Y(memwrite) );
	BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(aluout_0__RAW), .Y(aluout[0]) );
	BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(aluout_1__RAW), .Y(aluout[1]) );
	BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(aluout_2__RAW), .Y(aluout[2]) );
	BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(aluout_3__RAW), .Y(aluout[3]) );
	BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(aluout_4__RAW), .Y(aluout[4]) );
	BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(aluout_5__RAW), .Y(aluout[5]) );
	BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(aluout_6__RAW), .Y(aluout[6]) );
	BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(aluout_7__RAW), .Y(aluout[7]) );
	BUFX2 BUFX2_42 ( .gnd(gnd), .vdd(vdd), .A(aluout_8__RAW), .Y(aluout[8]) );
	BUFX2 BUFX2_43 ( .gnd(gnd), .vdd(vdd), .A(aluout_9__RAW), .Y(aluout[9]) );
	BUFX2 BUFX2_44 ( .gnd(gnd), .vdd(vdd), .A(aluout_10__RAW), .Y(aluout[10]) );
	BUFX2 BUFX2_45 ( .gnd(gnd), .vdd(vdd), .A(aluout_11__RAW), .Y(aluout[11]) );
	BUFX2 BUFX2_46 ( .gnd(gnd), .vdd(vdd), .A(aluout_12__RAW), .Y(aluout[12]) );
	BUFX2 BUFX2_47 ( .gnd(gnd), .vdd(vdd), .A(aluout_13__RAW), .Y(aluout[13]) );
	BUFX2 BUFX2_48 ( .gnd(gnd), .vdd(vdd), .A(aluout_14__RAW), .Y(aluout[14]) );
	BUFX2 BUFX2_49 ( .gnd(gnd), .vdd(vdd), .A(aluout_15__RAW), .Y(aluout[15]) );
	BUFX2 BUFX2_50 ( .gnd(gnd), .vdd(vdd), .A(aluout_16__RAW), .Y(aluout[16]) );
	BUFX2 BUFX2_51 ( .gnd(gnd), .vdd(vdd), .A(aluout_17__RAW), .Y(aluout[17]) );
	BUFX2 BUFX2_52 ( .gnd(gnd), .vdd(vdd), .A(aluout_18__RAW), .Y(aluout[18]) );
	BUFX2 BUFX2_53 ( .gnd(gnd), .vdd(vdd), .A(aluout_19__RAW), .Y(aluout[19]) );
	BUFX2 BUFX2_54 ( .gnd(gnd), .vdd(vdd), .A(aluout_20__RAW), .Y(aluout[20]) );
	BUFX2 BUFX2_55 ( .gnd(gnd), .vdd(vdd), .A(aluout_21__RAW), .Y(aluout[21]) );
	BUFX2 BUFX2_56 ( .gnd(gnd), .vdd(vdd), .A(aluout_22__RAW), .Y(aluout[22]) );
	BUFX2 BUFX2_57 ( .gnd(gnd), .vdd(vdd), .A(aluout_23__RAW), .Y(aluout[23]) );
	BUFX2 BUFX2_58 ( .gnd(gnd), .vdd(vdd), .A(aluout_24__RAW), .Y(aluout[24]) );
	BUFX2 BUFX2_59 ( .gnd(gnd), .vdd(vdd), .A(aluout_25__RAW), .Y(aluout[25]) );
	BUFX2 BUFX2_60 ( .gnd(gnd), .vdd(vdd), .A(aluout_26__RAW), .Y(aluout[26]) );
	BUFX2 BUFX2_61 ( .gnd(gnd), .vdd(vdd), .A(aluout_27__RAW), .Y(aluout[27]) );
	BUFX2 BUFX2_62 ( .gnd(gnd), .vdd(vdd), .A(aluout_28__RAW), .Y(aluout[28]) );
	BUFX2 BUFX2_63 ( .gnd(gnd), .vdd(vdd), .A(aluout_29__RAW), .Y(aluout[29]) );
	BUFX2 BUFX2_64 ( .gnd(gnd), .vdd(vdd), .A(aluout_30__RAW), .Y(aluout[30]) );
	BUFX2 BUFX2_65 ( .gnd(gnd), .vdd(vdd), .A(aluout_31__RAW), .Y(aluout[31]) );
	BUFX2 BUFX2_66 ( .gnd(gnd), .vdd(vdd), .A(writedata_0__RAW), .Y(writedata[0]) );
	BUFX2 BUFX2_67 ( .gnd(gnd), .vdd(vdd), .A(writedata_1__RAW), .Y(writedata[1]) );
	BUFX2 BUFX2_68 ( .gnd(gnd), .vdd(vdd), .A(writedata_2__RAW), .Y(writedata[2]) );
	BUFX2 BUFX2_69 ( .gnd(gnd), .vdd(vdd), .A(writedata_3__RAW), .Y(writedata[3]) );
	BUFX2 BUFX2_70 ( .gnd(gnd), .vdd(vdd), .A(writedata_4__RAW), .Y(writedata[4]) );
	BUFX2 BUFX2_71 ( .gnd(gnd), .vdd(vdd), .A(writedata_5__RAW), .Y(writedata[5]) );
	BUFX2 BUFX2_72 ( .gnd(gnd), .vdd(vdd), .A(writedata_6__RAW), .Y(writedata[6]) );
	BUFX2 BUFX2_73 ( .gnd(gnd), .vdd(vdd), .A(writedata_7__RAW), .Y(writedata[7]) );
	BUFX2 BUFX2_74 ( .gnd(gnd), .vdd(vdd), .A(writedata_8__RAW), .Y(writedata[8]) );
	BUFX2 BUFX2_75 ( .gnd(gnd), .vdd(vdd), .A(writedata_9__RAW), .Y(writedata[9]) );
	BUFX2 BUFX2_76 ( .gnd(gnd), .vdd(vdd), .A(writedata_10__RAW), .Y(writedata[10]) );
	BUFX2 BUFX2_77 ( .gnd(gnd), .vdd(vdd), .A(writedata_11__RAW), .Y(writedata[11]) );
	BUFX2 BUFX2_78 ( .gnd(gnd), .vdd(vdd), .A(writedata_12__RAW), .Y(writedata[12]) );
	BUFX2 BUFX2_79 ( .gnd(gnd), .vdd(vdd), .A(writedata_13__RAW), .Y(writedata[13]) );
	BUFX2 BUFX2_80 ( .gnd(gnd), .vdd(vdd), .A(writedata_14__RAW), .Y(writedata[14]) );
	BUFX2 BUFX2_81 ( .gnd(gnd), .vdd(vdd), .A(writedata_15__RAW), .Y(writedata[15]) );
	BUFX2 BUFX2_82 ( .gnd(gnd), .vdd(vdd), .A(writedata_16__RAW), .Y(writedata[16]) );
	BUFX2 BUFX2_83 ( .gnd(gnd), .vdd(vdd), .A(writedata_17__RAW), .Y(writedata[17]) );
	BUFX2 BUFX2_84 ( .gnd(gnd), .vdd(vdd), .A(writedata_18__RAW), .Y(writedata[18]) );
	BUFX2 BUFX2_85 ( .gnd(gnd), .vdd(vdd), .A(writedata_19__RAW), .Y(writedata[19]) );
	BUFX2 BUFX2_86 ( .gnd(gnd), .vdd(vdd), .A(writedata_20__RAW), .Y(writedata[20]) );
	BUFX2 BUFX2_87 ( .gnd(gnd), .vdd(vdd), .A(writedata_21__RAW), .Y(writedata[21]) );
	BUFX2 BUFX2_88 ( .gnd(gnd), .vdd(vdd), .A(writedata_22__RAW), .Y(writedata[22]) );
	BUFX2 BUFX2_89 ( .gnd(gnd), .vdd(vdd), .A(writedata_23__RAW), .Y(writedata[23]) );
	BUFX2 BUFX2_90 ( .gnd(gnd), .vdd(vdd), .A(writedata_24__RAW), .Y(writedata[24]) );
	BUFX2 BUFX2_91 ( .gnd(gnd), .vdd(vdd), .A(writedata_25__RAW), .Y(writedata[25]) );
	BUFX2 BUFX2_92 ( .gnd(gnd), .vdd(vdd), .A(writedata_26__RAW), .Y(writedata[26]) );
	BUFX2 BUFX2_93 ( .gnd(gnd), .vdd(vdd), .A(writedata_27__RAW), .Y(writedata[27]) );
	BUFX2 BUFX2_94 ( .gnd(gnd), .vdd(vdd), .A(writedata_28__RAW), .Y(writedata[28]) );
	BUFX2 BUFX2_95 ( .gnd(gnd), .vdd(vdd), .A(writedata_29__RAW), .Y(writedata[29]) );
	BUFX2 BUFX2_96 ( .gnd(gnd), .vdd(vdd), .A(writedata_30__RAW), .Y(writedata[30]) );
	BUFX2 BUFX2_97 ( .gnd(gnd), .vdd(vdd), .A(writedata_31__RAW), .Y(writedata[31]) );
	AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_0_), .B(zero), .Y(pcsrc) );
	INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(instr[2]), .Y(c.ad._abc_6357_n11_1) );
	AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n11_1), .B(instr[3]), .Y(c.ad._abc_6357_n12) );
	INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(instr[4]), .Y(c.ad._abc_6357_n13) );
	NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(instr[5]), .B(c.ad._abc_6357_n13), .Y(c.ad._abc_6357_n14) );
	INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(instr[0]), .Y(c.ad._abc_6357_n15) );
	NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(instr[1]), .B(c.ad._abc_6357_n15), .Y(c.ad._abc_6357_n16) );
	NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n14), .B(c.ad._abc_6357_n16), .Y(c.ad._abc_6357_n17) );
	NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n12), .B(c.ad._abc_6357_n17), .Y(c.ad._abc_6357_n18) );
	NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(instr[3]), .B(c.ad._abc_6357_n11_1), .Y(c.ad._abc_6357_n19) );
	INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(instr[1]), .Y(c.ad._abc_6357_n20) );
	NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(instr[0]), .B(c.ad._abc_6357_n20), .Y(c.ad._abc_6357_n21) );
	NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n14), .B(c.ad._abc_6357_n21), .Y(c.ad._abc_6357_n22) );
	NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n19), .B(c.ad._abc_6357_n22), .Y(c.ad._abc_6357_n23) );
	NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n18), .B(c.ad._abc_6357_n23), .Y(c.ad._abc_6357_n24) );
	AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n24), .B(c.aluop_1_), .Y(alucontrol_0_) );
	NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(instr[3]), .B(instr[2]), .Y(c.ad._abc_6357_n26_1) );
	NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n20), .B(c.ad._abc_6357_n15), .Y(c.ad._abc_6357_n27) );
	NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n14), .B(c.ad._abc_6357_n27), .Y(c.ad._abc_6357_n28) );
	NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n26_1), .B(c.ad._abc_6357_n28), .Y(c.ad._abc_6357_n29) );
	INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_1_), .Y(c.ad._abc_6357_n30) );
	NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(instr[0]), .B(c.ad._abc_6357_n20), .Y(c.ad._abc_6357_n31) );
	NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n11_1), .B(c.ad._abc_6357_n31), .Y(c.ad._abc_6357_n32) );
	NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n14), .B(c.ad._abc_6357_n32), .Y(c.ad._abc_6357_n33) );
	NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n30), .B(c.ad._abc_6357_n33), .Y(c.ad._abc_6357_n34) );
	NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n29), .B(c.ad._abc_6357_n34), .Y(alucontrol_1_) );
	NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_0_), .B(c.ad._abc_6357_n30), .Y(c.ad._abc_6357_n36) );
	NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_1_), .B(c.ad._abc_6357_n33), .Y(c.ad._abc_6357_n37) );
	NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(c.ad._abc_6357_n36), .B(c.ad._abc_6357_n37), .Y(alucontrol_2_) );
	INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(instr[29]), .Y(c.md._abc_6360_n13) );
	NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(instr[28]), .B(c.md._abc_6360_n13), .Y(c.md._abc_6360_n14) );
	NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(instr[27]), .B(instr[26]), .Y(c.md._abc_6360_n15) );
	NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(instr[31]), .B(instr[30]), .Y(c.md._abc_6360_n16) );
	NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n15), .B(c.md._abc_6360_n16), .Y(c.md._abc_6360_n17) );
	NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n14), .B(c.md._abc_6360_n17), .Y(c.aluop_0_) );
	NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(instr[29]), .B(instr[28]), .Y(c.md._abc_6360_n19) );
	INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n19), .Y(c.md._abc_6360_n20) );
	NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n20), .B(c.md._abc_6360_n17), .Y(c.aluop_1_) );
	INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(instr[26]), .Y(c.md._abc_6360_n22) );
	NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(instr[27]), .B(c.md._abc_6360_n22), .Y(c.md._abc_6360_n23) );
	NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n16), .B(c.md._abc_6360_n19), .Y(c.md._abc_6360_n24) );
	NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n23), .B(c.md._abc_6360_n24), .Y(c.md.controls_2_) );
	INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(instr[30]), .Y(c.md._abc_6360_n26) );
	NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(instr[31]), .B(c.md._abc_6360_n26), .Y(c.md._abc_6360_n27_1) );
	NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(instr[27]), .B(instr[26]), .Y(c.md._abc_6360_n28) );
	INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n28), .Y(c.md._abc_6360_n29) );
	NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n19), .B(c.md._abc_6360_n29), .Y(c.md._abc_6360_n30) );
	NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n27_1), .B(c.md._abc_6360_n30), .Y(c.md.controls_3_) );
	NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(instr[28]), .B(c.md._abc_6360_n13), .Y(c.md._abc_6360_n32) );
	NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n28), .B(c.md._abc_6360_n27_1), .Y(c.md._abc_6360_n33) );
	NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n32), .B(c.md._abc_6360_n33), .Y(c.md._abc_6360_n34) );
	INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n34), .Y(memwrite_RAW) );
	INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .Y(c.md._abc_6360_n36) );
	AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n15), .B(c.md._abc_6360_n16), .Y(c.md._abc_6360_n37) );
	NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n32), .B(c.md._abc_6360_n37), .Y(c.md._abc_6360_n38) );
	AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n34), .B(c.md._abc_6360_n38), .Y(c.md._abc_6360_n39) );
	NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n36), .B(c.md._abc_6360_n39), .Y(alusrc) );
	NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_1_), .B(c.md.controls_3_), .Y(c.md._abc_6360_n41) );
	NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(c.md._abc_6360_n38), .B(c.md._abc_6360_n41), .Y(c.md.controls_8_) );
	NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_1_), .B(alucontrol_0_), .Y(dp.alu._abc_6356_n100) );
	INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_1_), .Y(dp.alu._abc_6356_n101) );
	NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_0_), .B(dp.alu._abc_6356_n101), .Y(dp.alu._abc_6356_n102) );
	NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_0_), .B(dp.alu._abc_6356_n101), .Y(dp.alu._abc_6356_n103_1) );
	INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .Y(dp.alu._abc_6356_n104) );
	NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n102), .B(dp.alu._abc_6356_n104), .Y(dp.alu._abc_6356_n105) );
	NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n100), .B(dp.alu._abc_6356_n105), .Y(dp.alu._abc_6356_n106) );
	XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_28_), .Y(dp.alu._abc_6356_n107) );
	NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_28_), .B(dp.alu._abc_6356_n107), .Y(dp.alu._abc_6356_n108) );
	XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n107), .B(dp.srca_28_), .Y(dp.alu._abc_6356_n109) );
	XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_27_), .Y(dp.alu._abc_6356_n110_1) );
	NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_27_), .B(dp.alu._abc_6356_n110_1), .Y(dp.alu._abc_6356_n111) );
	XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n110_1), .B(dp.srca_27_), .Y(dp.alu._abc_6356_n112) );
	XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_26_), .Y(dp.alu._abc_6356_n113) );
	NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_26_), .B(dp.alu._abc_6356_n113), .Y(dp.alu._abc_6356_n114) );
	XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n113), .B(dp.srca_26_), .Y(dp.alu._abc_6356_n115) );
	XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_25_), .Y(dp.alu._abc_6356_n116) );
	NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_25_), .B(dp.alu._abc_6356_n116), .Y(dp.alu._abc_6356_n117_1) );
	XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n116), .B(dp.srca_25_), .Y(dp.alu._abc_6356_n118) );
	XOR2X1 XOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_24_), .Y(dp.alu._abc_6356_n119) );
	NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_24_), .B(dp.alu._abc_6356_n119), .Y(dp.alu._abc_6356_n120) );
	XOR2X1 XOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n119), .B(dp.srca_24_), .Y(dp.alu._abc_6356_n121) );
	XOR2X1 XOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_23_), .Y(dp.alu._abc_6356_n122) );
	NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_23_), .B(dp.alu._abc_6356_n122), .Y(dp.alu._abc_6356_n123) );
	XOR2X1 XOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n122), .B(dp.srca_23_), .Y(dp.alu._abc_6356_n124_1) );
	XOR2X1 XOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_22_), .Y(dp.alu._abc_6356_n125) );
	NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_22_), .B(dp.alu._abc_6356_n125), .Y(dp.alu._abc_6356_n126) );
	XOR2X1 XOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n125), .B(dp.srca_22_), .Y(dp.alu._abc_6356_n127) );
	XOR2X1 XOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_21_), .Y(dp.alu._abc_6356_n128) );
	NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_21_), .B(dp.alu._abc_6356_n128), .Y(dp.alu._abc_6356_n129) );
	XOR2X1 XOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n128), .B(dp.srca_21_), .Y(dp.alu._abc_6356_n130) );
	XOR2X1 XOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_20_), .Y(dp.alu._abc_6356_n131_1) );
	NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_20_), .B(dp.alu._abc_6356_n131_1), .Y(dp.alu._abc_6356_n132) );
	XOR2X1 XOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n131_1), .B(dp.srca_20_), .Y(dp.alu._abc_6356_n133) );
	XOR2X1 XOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_19_), .Y(dp.alu._abc_6356_n134) );
	NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_19_), .B(dp.alu._abc_6356_n134), .Y(dp.alu._abc_6356_n135) );
	XOR2X1 XOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n134), .B(dp.srca_19_), .Y(dp.alu._abc_6356_n136) );
	XOR2X1 XOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_18_), .Y(dp.alu._abc_6356_n137) );
	NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_18_), .B(dp.alu._abc_6356_n137), .Y(dp.alu._abc_6356_n138_1) );
	XOR2X1 XOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n137), .B(dp.srca_18_), .Y(dp.alu._abc_6356_n139) );
	XOR2X1 XOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_17_), .Y(dp.alu._abc_6356_n140) );
	NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_17_), .B(dp.alu._abc_6356_n140), .Y(dp.alu._abc_6356_n141) );
	XOR2X1 XOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n140), .B(dp.srca_17_), .Y(dp.alu._abc_6356_n142) );
	XOR2X1 XOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_16_), .Y(dp.alu._abc_6356_n143) );
	NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_16_), .B(dp.alu._abc_6356_n143), .Y(dp.alu._abc_6356_n144) );
	XOR2X1 XOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n143), .B(dp.srca_16_), .Y(dp.alu._abc_6356_n145_1) );
	XOR2X1 XOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_15_), .Y(dp.alu._abc_6356_n146) );
	NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_15_), .B(dp.alu._abc_6356_n146), .Y(dp.alu._abc_6356_n147) );
	XOR2X1 XOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n146), .B(dp.srca_15_), .Y(dp.alu._abc_6356_n148) );
	XOR2X1 XOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_14_), .Y(dp.alu._abc_6356_n149) );
	NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_14_), .B(dp.alu._abc_6356_n149), .Y(dp.alu._abc_6356_n150) );
	XOR2X1 XOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n149), .B(dp.srca_14_), .Y(dp.alu._abc_6356_n151) );
	XOR2X1 XOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_13_), .Y(dp.alu._abc_6356_n152_1) );
	NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_13_), .B(dp.alu._abc_6356_n152_1), .Y(dp.alu._abc_6356_n153) );
	XOR2X1 XOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n152_1), .B(dp.srca_13_), .Y(dp.alu._abc_6356_n154) );
	XOR2X1 XOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_12_), .Y(dp.alu._abc_6356_n155) );
	NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_12_), .B(dp.alu._abc_6356_n155), .Y(dp.alu._abc_6356_n156) );
	XOR2X1 XOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n155), .B(dp.srca_12_), .Y(dp.alu._abc_6356_n157) );
	XOR2X1 XOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_11_), .Y(dp.alu._abc_6356_n158) );
	NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_11_), .B(dp.alu._abc_6356_n158), .Y(dp.alu._abc_6356_n159_1) );
	XOR2X1 XOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n158), .B(dp.srca_11_), .Y(dp.alu._abc_6356_n160) );
	XOR2X1 XOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_10_), .Y(dp.alu._abc_6356_n161) );
	NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_10_), .B(dp.alu._abc_6356_n161), .Y(dp.alu._abc_6356_n162) );
	XOR2X1 XOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n161), .B(dp.srca_10_), .Y(dp.alu._abc_6356_n163) );
	XOR2X1 XOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_9_), .Y(dp.alu._abc_6356_n164) );
	NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_9_), .B(dp.alu._abc_6356_n164), .Y(dp.alu._abc_6356_n165) );
	XOR2X1 XOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n164), .B(dp.srca_9_), .Y(dp.alu._abc_6356_n166_1) );
	XOR2X1 XOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_8_), .Y(dp.alu._abc_6356_n167) );
	NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_8_), .B(dp.alu._abc_6356_n167), .Y(dp.alu._abc_6356_n168) );
	XOR2X1 XOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n167), .B(dp.srca_8_), .Y(dp.alu._abc_6356_n169) );
	XOR2X1 XOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_7_), .Y(dp.alu._abc_6356_n170_1) );
	NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_7_), .B(dp.alu._abc_6356_n170_1), .Y(dp.alu._abc_6356_n171) );
	XOR2X1 XOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n170_1), .B(dp.srca_7_), .Y(dp.alu._abc_6356_n172) );
	XOR2X1 XOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_6_), .Y(dp.alu._abc_6356_n173) );
	NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_6_), .B(dp.alu._abc_6356_n173), .Y(dp.alu._abc_6356_n174) );
	XOR2X1 XOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n173), .B(dp.srca_6_), .Y(dp.alu._abc_6356_n175) );
	XOR2X1 XOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_5_), .Y(dp.alu._abc_6356_n176) );
	NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_5_), .B(dp.alu._abc_6356_n176), .Y(dp.alu._abc_6356_n177_1) );
	XOR2X1 XOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n176), .B(dp.srca_5_), .Y(dp.alu._abc_6356_n178) );
	XOR2X1 XOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_4_), .Y(dp.alu._abc_6356_n179) );
	NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_4_), .B(dp.alu._abc_6356_n179), .Y(dp.alu._abc_6356_n180) );
	XOR2X1 XOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n179), .B(dp.srca_4_), .Y(dp.alu._abc_6356_n181) );
	XOR2X1 XOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_3_), .Y(dp.alu._abc_6356_n182) );
	NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_3_), .B(dp.alu._abc_6356_n182), .Y(dp.alu._abc_6356_n183) );
	XOR2X1 XOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n182), .B(dp.srca_3_), .Y(dp.alu._abc_6356_n184_1) );
	XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_2_), .Y(dp.alu._abc_6356_n185) );
	INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n185), .Y(dp.alu._abc_6356_n186) );
	NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_2_), .B(dp.alu._abc_6356_n186), .Y(dp.alu._abc_6356_n187) );
	XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n185), .B(dp.srca_2_), .Y(dp.alu._abc_6356_n188) );
	NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_1_), .Y(dp.alu._abc_6356_n189) );
	AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_1_), .Y(dp.alu._abc_6356_n190) );
	NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n189), .B(dp.alu._abc_6356_n190), .Y(dp.alu._abc_6356_n191_1) );
	NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_1_), .B(dp.alu._abc_6356_n191_1), .Y(dp.alu._abc_6356_n192) );
	NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_0_), .Y(dp.alu._abc_6356_n193) );
	NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_0_), .Y(dp.alu._abc_6356_n194) );
	NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_0_), .B(dp.alu._abc_6356_n194), .Y(dp.alu._abc_6356_n195) );
	NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n193), .B(dp.alu._abc_6356_n195), .Y(dp.alu._abc_6356_n196) );
	INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_1_), .Y(dp.alu._abc_6356_n197) );
	NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n197), .B(dp.alu._abc_6356_n191_1), .Y(dp.alu._abc_6356_n198_1) );
	XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_1_), .Y(dp.alu._abc_6356_n199) );
	NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_1_), .B(dp.alu._abc_6356_n199), .Y(dp.alu._abc_6356_n200) );
	NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n198_1), .B(dp.alu._abc_6356_n200), .Y(dp.alu._abc_6356_n201) );
	NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n196), .B(dp.alu._abc_6356_n201), .Y(dp.alu._abc_6356_n202) );
	NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n192), .B(dp.alu._abc_6356_n202), .Y(dp.alu._abc_6356_n203) );
	NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n188), .B(dp.alu._abc_6356_n203), .Y(dp.alu._abc_6356_n204) );
	NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n187), .B(dp.alu._abc_6356_n204), .Y(dp.alu._abc_6356_n205_1) );
	NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n184_1), .B(dp.alu._abc_6356_n205_1), .Y(dp.alu._abc_6356_n206) );
	NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n183), .B(dp.alu._abc_6356_n206), .Y(dp.alu._abc_6356_n207) );
	NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n181), .B(dp.alu._abc_6356_n207), .Y(dp.alu._abc_6356_n208) );
	NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n180), .B(dp.alu._abc_6356_n208), .Y(dp.alu._abc_6356_n209) );
	NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n178), .B(dp.alu._abc_6356_n209), .Y(dp.alu._abc_6356_n210) );
	NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n177_1), .B(dp.alu._abc_6356_n210), .Y(dp.alu._abc_6356_n211) );
	NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n175), .B(dp.alu._abc_6356_n211), .Y(dp.alu._abc_6356_n212_1) );
	NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n174), .B(dp.alu._abc_6356_n212_1), .Y(dp.alu._abc_6356_n213) );
	NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n172), .B(dp.alu._abc_6356_n213), .Y(dp.alu._abc_6356_n214) );
	NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n171), .B(dp.alu._abc_6356_n214), .Y(dp.alu._abc_6356_n215) );
	NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n169), .B(dp.alu._abc_6356_n215), .Y(dp.alu._abc_6356_n216) );
	NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n168), .B(dp.alu._abc_6356_n216), .Y(dp.alu._abc_6356_n217) );
	NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n166_1), .B(dp.alu._abc_6356_n217), .Y(dp.alu._abc_6356_n218_1) );
	NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n165), .B(dp.alu._abc_6356_n218_1), .Y(dp.alu._abc_6356_n219) );
	NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n163), .B(dp.alu._abc_6356_n219), .Y(dp.alu._abc_6356_n220) );
	NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n162), .B(dp.alu._abc_6356_n220), .Y(dp.alu._abc_6356_n221) );
	NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n160), .B(dp.alu._abc_6356_n221), .Y(dp.alu._abc_6356_n222) );
	NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n159_1), .B(dp.alu._abc_6356_n222), .Y(dp.alu._abc_6356_n223) );
	NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n157), .B(dp.alu._abc_6356_n223), .Y(dp.alu._abc_6356_n224) );
	NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n156), .B(dp.alu._abc_6356_n224), .Y(dp.alu._abc_6356_n225) );
	NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n154), .B(dp.alu._abc_6356_n225), .Y(dp.alu._abc_6356_n226) );
	NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n153), .B(dp.alu._abc_6356_n226), .Y(dp.alu._abc_6356_n227) );
	NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n151), .B(dp.alu._abc_6356_n227), .Y(dp.alu._abc_6356_n228) );
	NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n150), .B(dp.alu._abc_6356_n228), .Y(dp.alu._abc_6356_n229) );
	NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n148), .B(dp.alu._abc_6356_n229), .Y(dp.alu._abc_6356_n230) );
	NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n147), .B(dp.alu._abc_6356_n230), .Y(dp.alu._abc_6356_n231) );
	NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n145_1), .B(dp.alu._abc_6356_n231), .Y(dp.alu._abc_6356_n232) );
	NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n144), .B(dp.alu._abc_6356_n232), .Y(dp.alu._abc_6356_n233) );
	NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n142), .B(dp.alu._abc_6356_n233), .Y(dp.alu._abc_6356_n234) );
	NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n141), .B(dp.alu._abc_6356_n234), .Y(dp.alu._abc_6356_n235) );
	NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n139), .B(dp.alu._abc_6356_n235), .Y(dp.alu._abc_6356_n236) );
	NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n138_1), .B(dp.alu._abc_6356_n236), .Y(dp.alu._abc_6356_n237) );
	NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n136), .B(dp.alu._abc_6356_n237), .Y(dp.alu._abc_6356_n238) );
	NAND2X1 NAND2X1_97 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n135), .B(dp.alu._abc_6356_n238), .Y(dp.alu._abc_6356_n239) );
	NAND2X1 NAND2X1_98 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n133), .B(dp.alu._abc_6356_n239), .Y(dp.alu._abc_6356_n240) );
	NAND2X1 NAND2X1_99 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n132), .B(dp.alu._abc_6356_n240), .Y(dp.alu._abc_6356_n241) );
	NAND2X1 NAND2X1_100 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n130), .B(dp.alu._abc_6356_n241), .Y(dp.alu._abc_6356_n242) );
	NAND2X1 NAND2X1_101 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n129), .B(dp.alu._abc_6356_n242), .Y(dp.alu._abc_6356_n243) );
	NAND2X1 NAND2X1_102 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n127), .B(dp.alu._abc_6356_n243), .Y(dp.alu._abc_6356_n244) );
	NAND2X1 NAND2X1_103 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n126), .B(dp.alu._abc_6356_n244), .Y(dp.alu._abc_6356_n245) );
	NAND2X1 NAND2X1_104 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n124_1), .B(dp.alu._abc_6356_n245), .Y(dp.alu._abc_6356_n246) );
	NAND2X1 NAND2X1_105 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n123), .B(dp.alu._abc_6356_n246), .Y(dp.alu._abc_6356_n247) );
	NAND2X1 NAND2X1_106 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n121), .B(dp.alu._abc_6356_n247), .Y(dp.alu._abc_6356_n248) );
	NAND2X1 NAND2X1_107 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n120), .B(dp.alu._abc_6356_n248), .Y(dp.alu._abc_6356_n249) );
	NAND2X1 NAND2X1_108 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n118), .B(dp.alu._abc_6356_n249), .Y(dp.alu._abc_6356_n250) );
	NAND2X1 NAND2X1_109 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n117_1), .B(dp.alu._abc_6356_n250), .Y(dp.alu._abc_6356_n251) );
	NAND2X1 NAND2X1_110 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n115), .B(dp.alu._abc_6356_n251), .Y(dp.alu._abc_6356_n252) );
	NAND2X1 NAND2X1_111 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n114), .B(dp.alu._abc_6356_n252), .Y(dp.alu._abc_6356_n253) );
	NAND2X1 NAND2X1_112 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n112), .B(dp.alu._abc_6356_n253), .Y(dp.alu._abc_6356_n254) );
	NAND2X1 NAND2X1_113 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n111), .B(dp.alu._abc_6356_n254), .Y(dp.alu._abc_6356_n255) );
	NAND2X1 NAND2X1_114 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n109), .B(dp.alu._abc_6356_n255), .Y(dp.alu._abc_6356_n256) );
	NAND2X1 NAND2X1_115 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n108), .B(dp.alu._abc_6356_n256), .Y(dp.alu._abc_6356_n257) );
	XOR2X1 XOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_29_), .Y(dp.alu._abc_6356_n258) );
	XOR2X1 XOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n258), .B(dp.srca_29_), .Y(dp.alu._abc_6356_n259) );
	XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n257), .B(dp.alu._abc_6356_n259), .Y(dp.alu._abc_6356_n260) );
	XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n255), .B(dp.alu._abc_6356_n109), .Y(dp.alu._abc_6356_n261) );
	XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n253), .B(dp.alu._abc_6356_n112), .Y(dp.alu._abc_6356_n262) );
	XOR2X1 XOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n251), .B(dp.alu._abc_6356_n115), .Y(dp.alu._abc_6356_n263) );
	XOR2X1 XOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n247), .B(dp.alu._abc_6356_n121), .Y(dp.alu._abc_6356_n264) );
	XOR2X1 XOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n243), .B(dp.alu._abc_6356_n127), .Y(dp.alu._abc_6356_n265) );
	XOR2X1 XOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n239), .B(dp.alu._abc_6356_n133), .Y(dp.alu._abc_6356_n266) );
	XOR2X1 XOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n235), .B(dp.alu._abc_6356_n139), .Y(dp.alu._abc_6356_n267) );
	XOR2X1 XOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n231), .B(dp.alu._abc_6356_n145_1), .Y(dp.alu._abc_6356_n268) );
	XOR2X1 XOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n227), .B(dp.alu._abc_6356_n151), .Y(dp.alu._abc_6356_n269) );
	XOR2X1 XOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n223), .B(dp.alu._abc_6356_n157), .Y(dp.alu._abc_6356_n270) );
	XOR2X1 XOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n219), .B(dp.alu._abc_6356_n163), .Y(dp.alu._abc_6356_n271) );
	XOR2X1 XOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n215), .B(dp.alu._abc_6356_n169), .Y(dp.alu._abc_6356_n272) );
	XOR2X1 XOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n205_1), .B(dp.alu._abc_6356_n184_1), .Y(dp.alu._abc_6356_n273) );
	INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .Y(dp.alu._abc_6356_n274) );
	NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_0_), .B(dp.srcb_0_), .Y(dp.alu._abc_6356_n275) );
	NAND2X1 NAND2X1_116 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_0_), .B(dp.srcb_0_), .Y(dp.alu._abc_6356_n276) );
	INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n276), .Y(dp.alu._abc_6356_n277) );
	NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n275), .B(dp.alu._abc_6356_n277), .Y(dp.alu._abc_6356_n278) );
	NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n274), .B(dp.alu._abc_6356_n278), .Y(dp.alu._abc_6356_n279) );
	XOR2X1 XOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n201), .B(dp.alu._abc_6356_n196), .Y(dp.alu._abc_6356_n280) );
	NAND2X1 NAND2X1_117 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n279), .B(dp.alu._abc_6356_n280), .Y(dp.alu._abc_6356_n281) );
	XOR2X1 XOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n203), .B(dp.alu._abc_6356_n188), .Y(dp.alu._abc_6356_n282) );
	INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n282), .Y(dp.alu._abc_6356_n283) );
	NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n281), .B(dp.alu._abc_6356_n283), .Y(dp.alu._abc_6356_n284) );
	NAND2X1 NAND2X1_118 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n273), .B(dp.alu._abc_6356_n284), .Y(dp.alu._abc_6356_n285) );
	INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n285), .Y(dp.alu._abc_6356_n286) );
	XOR2X1 XOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n207), .B(dp.alu._abc_6356_n181), .Y(dp.alu._abc_6356_n287) );
	NAND2X1 NAND2X1_119 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n286), .B(dp.alu._abc_6356_n287), .Y(dp.alu._abc_6356_n288) );
	INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n288), .Y(dp.alu._abc_6356_n289) );
	XOR2X1 XOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n209), .B(dp.alu._abc_6356_n178), .Y(dp.alu._abc_6356_n290) );
	NAND2X1 NAND2X1_120 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n289), .B(dp.alu._abc_6356_n290), .Y(dp.alu._abc_6356_n291) );
	INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n291), .Y(dp.alu._abc_6356_n292) );
	XOR2X1 XOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n211), .B(dp.alu._abc_6356_n175), .Y(dp.alu._abc_6356_n293) );
	NAND2X1 NAND2X1_121 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n292), .B(dp.alu._abc_6356_n293), .Y(dp.alu._abc_6356_n294) );
	XOR2X1 XOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n213), .B(dp.alu._abc_6356_n172), .Y(dp.alu._abc_6356_n295) );
	INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n295), .Y(dp.alu._abc_6356_n296) );
	NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n294), .B(dp.alu._abc_6356_n296), .Y(dp.alu._abc_6356_n297) );
	NAND2X1 NAND2X1_122 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n272), .B(dp.alu._abc_6356_n297), .Y(dp.alu._abc_6356_n298) );
	XOR2X1 XOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n217), .B(dp.alu._abc_6356_n166_1), .Y(dp.alu._abc_6356_n299) );
	INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n299), .Y(dp.alu._abc_6356_n300) );
	NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n298), .B(dp.alu._abc_6356_n300), .Y(dp.alu._abc_6356_n301) );
	NAND2X1 NAND2X1_123 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n271), .B(dp.alu._abc_6356_n301), .Y(dp.alu._abc_6356_n302) );
	XOR2X1 XOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n221), .B(dp.alu._abc_6356_n160), .Y(dp.alu._abc_6356_n303) );
	INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n303), .Y(dp.alu._abc_6356_n304) );
	NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n302), .B(dp.alu._abc_6356_n304), .Y(dp.alu._abc_6356_n305) );
	NAND2X1 NAND2X1_124 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n270), .B(dp.alu._abc_6356_n305), .Y(dp.alu._abc_6356_n306) );
	XOR2X1 XOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n225), .B(dp.alu._abc_6356_n154), .Y(dp.alu._abc_6356_n307) );
	INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n307), .Y(dp.alu._abc_6356_n308) );
	NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n306), .B(dp.alu._abc_6356_n308), .Y(dp.alu._abc_6356_n309) );
	NAND2X1 NAND2X1_125 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n269), .B(dp.alu._abc_6356_n309), .Y(dp.alu._abc_6356_n310) );
	XOR2X1 XOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n229), .B(dp.alu._abc_6356_n148), .Y(dp.alu._abc_6356_n311) );
	INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n311), .Y(dp.alu._abc_6356_n312) );
	NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n310), .B(dp.alu._abc_6356_n312), .Y(dp.alu._abc_6356_n313) );
	NAND2X1 NAND2X1_126 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n268), .B(dp.alu._abc_6356_n313), .Y(dp.alu._abc_6356_n314) );
	XOR2X1 XOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n233), .B(dp.alu._abc_6356_n142), .Y(dp.alu._abc_6356_n315) );
	INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n315), .Y(dp.alu._abc_6356_n316) );
	NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n314), .B(dp.alu._abc_6356_n316), .Y(dp.alu._abc_6356_n317) );
	NAND2X1 NAND2X1_127 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n267), .B(dp.alu._abc_6356_n317), .Y(dp.alu._abc_6356_n318) );
	XOR2X1 XOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n237), .B(dp.alu._abc_6356_n136), .Y(dp.alu._abc_6356_n319) );
	INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n319), .Y(dp.alu._abc_6356_n320) );
	NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n318), .B(dp.alu._abc_6356_n320), .Y(dp.alu._abc_6356_n321) );
	NAND2X1 NAND2X1_128 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n266), .B(dp.alu._abc_6356_n321), .Y(dp.alu._abc_6356_n322) );
	XOR2X1 XOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n241), .B(dp.alu._abc_6356_n130), .Y(dp.alu._abc_6356_n323) );
	INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n323), .Y(dp.alu._abc_6356_n324) );
	NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n322), .B(dp.alu._abc_6356_n324), .Y(dp.alu._abc_6356_n325) );
	NAND2X1 NAND2X1_129 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n265), .B(dp.alu._abc_6356_n325), .Y(dp.alu._abc_6356_n326) );
	XOR2X1 XOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n245), .B(dp.alu._abc_6356_n124_1), .Y(dp.alu._abc_6356_n327) );
	INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n327), .Y(dp.alu._abc_6356_n328) );
	NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n326), .B(dp.alu._abc_6356_n328), .Y(dp.alu._abc_6356_n329) );
	NAND2X1 NAND2X1_130 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n264), .B(dp.alu._abc_6356_n329), .Y(dp.alu._abc_6356_n330) );
	XOR2X1 XOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n249), .B(dp.alu._abc_6356_n118), .Y(dp.alu._abc_6356_n331) );
	INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n331), .Y(dp.alu._abc_6356_n332) );
	NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n330), .B(dp.alu._abc_6356_n332), .Y(dp.alu._abc_6356_n333) );
	NAND2X1 NAND2X1_131 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n263), .B(dp.alu._abc_6356_n333), .Y(dp.alu._abc_6356_n334) );
	OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n262), .B(dp.alu._abc_6356_n334), .Y(dp.alu._abc_6356_n335) );
	OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n261), .B(dp.alu._abc_6356_n335), .Y(dp.alu._abc_6356_n336) );
	OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n260), .B(dp.alu._abc_6356_n336), .Y(dp.alu._abc_6356_n337) );
	NAND2X1 NAND2X1_132 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_29_), .B(dp.alu._abc_6356_n258), .Y(dp.alu._abc_6356_n338) );
	NAND2X1 NAND2X1_133 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n259), .B(dp.alu._abc_6356_n257), .Y(dp.alu._abc_6356_n339) );
	NAND2X1 NAND2X1_134 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n338), .B(dp.alu._abc_6356_n339), .Y(dp.alu._abc_6356_n340) );
	XOR2X1 XOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_2_), .B(dp.srcb_30_), .Y(dp.alu._abc_6356_n341) );
	XOR2X1 XOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n341), .B(dp.srca_30_), .Y(dp.alu._abc_6356_n342) );
	XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n340), .B(dp.alu._abc_6356_n342), .Y(dp.alu._abc_6356_n343) );
	NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n337), .B(dp.alu._abc_6356_n343), .Y(dp.alu._abc_6356_n344) );
	NAND2X1 NAND2X1_135 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_30_), .B(dp.alu._abc_6356_n341), .Y(dp.alu._abc_6356_n345) );
	NAND2X1 NAND2X1_136 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n342), .B(dp.alu._abc_6356_n340), .Y(dp.alu._abc_6356_n346) );
	NAND2X1 NAND2X1_137 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n345), .B(dp.alu._abc_6356_n346), .Y(dp.alu._abc_6356_n347) );
	NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_31_), .B(dp.srcb_31_), .Y(dp.alu._abc_6356_n348) );
	NAND2X1 NAND2X1_138 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_31_), .B(dp.srcb_31_), .Y(dp.alu._abc_6356_n349) );
	INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n349), .Y(dp.alu._abc_6356_n350) );
	NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n348), .B(dp.alu._abc_6356_n350), .Y(dp.alu._abc_6356_n351) );
	XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n351), .B(alucontrol_2_), .Y(dp.alu._abc_6356_n352) );
	INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n352), .Y(dp.alu._abc_6356_n353) );
	XNOR2X1 XNOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n347), .B(dp.alu._abc_6356_n353), .Y(dp.alu._abc_6356_n354) );
	NAND2X1 NAND2X1_139 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n344), .B(dp.alu._abc_6356_n354), .Y(dp.alu._abc_6356_n355) );
	OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n343), .B(dp.alu._abc_6356_n337), .Y(dp.alu._abc_6356_n356) );
	XNOR2X1 XNOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n347), .B(dp.alu._abc_6356_n352), .Y(dp.alu._abc_6356_n357) );
	NAND2X1 NAND2X1_140 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n356), .B(dp.alu._abc_6356_n357), .Y(dp.alu._abc_6356_n358) );
	NAND2X1 NAND2X1_141 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n355), .B(dp.alu._abc_6356_n358), .Y(dp.alu._abc_6356_n359) );
	NAND2X1 NAND2X1_142 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n106), .B(dp.alu._abc_6356_n359), .Y(dp.alu._abc_6356_n360) );
	NAND2X1 NAND2X1_143 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n278), .B(dp.alu._abc_6356_n105), .Y(dp.alu._abc_6356_n361) );
	NAND2X1 NAND2X1_144 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n101), .B(dp.alu._abc_6356_n277), .Y(dp.alu._abc_6356_n362) );
	AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n361), .B(dp.alu._abc_6356_n362), .Y(dp.alu._abc_6356_n363) );
	AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n360), .B(dp.alu._abc_6356_n363), .Y(dp.alu._abc_6356_n364) );
	INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n364), .Y(aluout_0__RAW) );
	AND2X2 AND2X2_9 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_1_), .B(dp.srcb_1_), .Y(dp.alu._abc_6356_n366) );
	AND2X2 AND2X2_10 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n366), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n367) );
	NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_1_), .B(dp.srcb_1_), .Y(dp.alu._abc_6356_n368) );
	NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n368), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n369) );
	NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n367), .B(dp.alu._abc_6356_n369), .Y(dp.alu._abc_6356_n370) );
	XOR2X1 XOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n280), .B(dp.alu._abc_6356_n279), .Y(dp.alu._abc_6356_n371) );
	NAND2X1 NAND2X1_145 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n371), .Y(dp.alu._abc_6356_n372) );
	NAND2X1 NAND2X1_146 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n370), .B(dp.alu._abc_6356_n372), .Y(aluout_1__RAW) );
	AND2X2 AND2X2_11 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_2_), .B(dp.srcb_2_), .Y(dp.alu._abc_6356_n374) );
	AND2X2 AND2X2_12 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n374), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n375) );
	NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_2_), .B(dp.srcb_2_), .Y(dp.alu._abc_6356_n376) );
	NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n376), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n377) );
	NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n375), .B(dp.alu._abc_6356_n377), .Y(dp.alu._abc_6356_n378) );
	NAND2X1 NAND2X1_147 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n281), .B(dp.alu._abc_6356_n283), .Y(dp.alu._abc_6356_n379) );
	NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n284), .Y(dp.alu._abc_6356_n380) );
	NAND2X1 NAND2X1_148 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n379), .B(dp.alu._abc_6356_n380), .Y(dp.alu._abc_6356_n381) );
	NAND2X1 NAND2X1_149 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n378), .B(dp.alu._abc_6356_n381), .Y(aluout_2__RAW) );
	AND2X2 AND2X2_13 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_3_), .B(dp.srcb_3_), .Y(dp.alu._abc_6356_n383) );
	AND2X2 AND2X2_14 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n383), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n384) );
	NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_3_), .B(dp.srcb_3_), .Y(dp.alu._abc_6356_n385) );
	NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n385), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n386) );
	NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n384), .B(dp.alu._abc_6356_n386), .Y(dp.alu._abc_6356_n387) );
	NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n273), .B(dp.alu._abc_6356_n284), .Y(dp.alu._abc_6356_n388) );
	NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n388), .B(dp.alu._abc_6356_n286), .Y(dp.alu._abc_6356_n389) );
	NAND2X1 NAND2X1_150 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n389), .Y(dp.alu._abc_6356_n390) );
	NAND2X1 NAND2X1_151 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n387), .B(dp.alu._abc_6356_n390), .Y(aluout_3__RAW) );
	AND2X2 AND2X2_15 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_4_), .B(dp.srcb_4_), .Y(dp.alu._abc_6356_n392) );
	AND2X2 AND2X2_16 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n392), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n393) );
	NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_4_), .B(dp.srcb_4_), .Y(dp.alu._abc_6356_n394) );
	NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n394), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n395) );
	NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n393), .B(dp.alu._abc_6356_n395), .Y(dp.alu._abc_6356_n396) );
	XNOR2X1 XNOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n287), .B(dp.alu._abc_6356_n285), .Y(dp.alu._abc_6356_n397) );
	NAND2X1 NAND2X1_152 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n397), .Y(dp.alu._abc_6356_n398) );
	NAND2X1 NAND2X1_153 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n396), .B(dp.alu._abc_6356_n398), .Y(aluout_4__RAW) );
	AND2X2 AND2X2_17 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_5_), .B(dp.srcb_5_), .Y(dp.alu._abc_6356_n400) );
	AND2X2 AND2X2_18 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n400), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n401) );
	NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_5_), .B(dp.srcb_5_), .Y(dp.alu._abc_6356_n402) );
	NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n402), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n403) );
	NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n401), .B(dp.alu._abc_6356_n403), .Y(dp.alu._abc_6356_n404) );
	NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n289), .B(dp.alu._abc_6356_n290), .Y(dp.alu._abc_6356_n405) );
	NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n405), .B(dp.alu._abc_6356_n292), .Y(dp.alu._abc_6356_n406) );
	NAND2X1 NAND2X1_154 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n406), .Y(dp.alu._abc_6356_n407) );
	NAND2X1 NAND2X1_155 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n404), .B(dp.alu._abc_6356_n407), .Y(aluout_5__RAW) );
	AND2X2 AND2X2_19 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_6_), .B(dp.srcb_6_), .Y(dp.alu._abc_6356_n409) );
	AND2X2 AND2X2_20 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n409), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n410) );
	NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_6_), .B(dp.srcb_6_), .Y(dp.alu._abc_6356_n411) );
	NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n411), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n412) );
	NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n410), .B(dp.alu._abc_6356_n412), .Y(dp.alu._abc_6356_n413) );
	XNOR2X1 XNOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n293), .B(dp.alu._abc_6356_n291), .Y(dp.alu._abc_6356_n414) );
	NAND2X1 NAND2X1_156 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n414), .Y(dp.alu._abc_6356_n415) );
	NAND2X1 NAND2X1_157 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n413), .B(dp.alu._abc_6356_n415), .Y(aluout_6__RAW) );
	AND2X2 AND2X2_21 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_7_), .B(dp.srcb_7_), .Y(dp.alu._abc_6356_n417) );
	AND2X2 AND2X2_22 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n417), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n418) );
	NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_7_), .B(dp.srcb_7_), .Y(dp.alu._abc_6356_n419) );
	NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n419), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n420) );
	NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n418), .B(dp.alu._abc_6356_n420), .Y(dp.alu._abc_6356_n421) );
	NAND2X1 NAND2X1_158 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n294), .B(dp.alu._abc_6356_n296), .Y(dp.alu._abc_6356_n422) );
	NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n297), .Y(dp.alu._abc_6356_n423) );
	NAND2X1 NAND2X1_159 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n422), .B(dp.alu._abc_6356_n423), .Y(dp.alu._abc_6356_n424) );
	NAND2X1 NAND2X1_160 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n421), .B(dp.alu._abc_6356_n424), .Y(aluout_7__RAW) );
	AND2X2 AND2X2_23 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_8_), .B(dp.srcb_8_), .Y(dp.alu._abc_6356_n426) );
	AND2X2 AND2X2_24 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n426), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n427) );
	NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_8_), .B(dp.srcb_8_), .Y(dp.alu._abc_6356_n428) );
	NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n428), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n429) );
	NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n427), .B(dp.alu._abc_6356_n429), .Y(dp.alu._abc_6356_n430) );
	NAND2X1 NAND2X1_161 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n298), .Y(dp.alu._abc_6356_n431) );
	NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n272), .B(dp.alu._abc_6356_n297), .Y(dp.alu._abc_6356_n432) );
	OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n431), .B(dp.alu._abc_6356_n432), .Y(dp.alu._abc_6356_n433) );
	NAND2X1 NAND2X1_162 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n430), .B(dp.alu._abc_6356_n433), .Y(aluout_8__RAW) );
	AND2X2 AND2X2_25 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_9_), .B(dp.srcb_9_), .Y(dp.alu._abc_6356_n435) );
	AND2X2 AND2X2_26 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n435), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n436) );
	NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_9_), .B(dp.srcb_9_), .Y(dp.alu._abc_6356_n437) );
	NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n437), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n438) );
	NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n436), .B(dp.alu._abc_6356_n438), .Y(dp.alu._abc_6356_n439) );
	NAND2X1 NAND2X1_163 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n298), .B(dp.alu._abc_6356_n300), .Y(dp.alu._abc_6356_n440) );
	NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n301), .Y(dp.alu._abc_6356_n441) );
	NAND2X1 NAND2X1_164 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n440), .B(dp.alu._abc_6356_n441), .Y(dp.alu._abc_6356_n442) );
	NAND2X1 NAND2X1_165 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n439), .B(dp.alu._abc_6356_n442), .Y(aluout_9__RAW) );
	AND2X2 AND2X2_27 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_10_), .B(dp.srcb_10_), .Y(dp.alu._abc_6356_n444) );
	AND2X2 AND2X2_28 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n444), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n445_1) );
	NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_10_), .B(dp.srcb_10_), .Y(dp.alu._abc_6356_n446) );
	NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n446), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n447) );
	NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n445_1), .B(dp.alu._abc_6356_n447), .Y(dp.alu._abc_6356_n448_1) );
	NAND2X1 NAND2X1_166 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n302), .Y(dp.alu._abc_6356_n449) );
	NOR2X1 NOR2X1_81 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n271), .B(dp.alu._abc_6356_n301), .Y(dp.alu._abc_6356_n450_1) );
	OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n449), .B(dp.alu._abc_6356_n450_1), .Y(dp.alu._abc_6356_n451_1) );
	NAND2X1 NAND2X1_167 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n448_1), .B(dp.alu._abc_6356_n451_1), .Y(aluout_10__RAW) );
	AND2X2 AND2X2_29 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_11_), .B(dp.srcb_11_), .Y(dp.alu._abc_6356_n453_1) );
	AND2X2 AND2X2_30 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n453_1), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n454_1) );
	NOR2X1 NOR2X1_82 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_11_), .B(dp.srcb_11_), .Y(dp.alu._abc_6356_n455_1) );
	NOR2X1 NOR2X1_83 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n455_1), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n456_1) );
	NOR2X1 NOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n454_1), .B(dp.alu._abc_6356_n456_1), .Y(dp.alu._abc_6356_n457_1) );
	NAND2X1 NAND2X1_168 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n302), .B(dp.alu._abc_6356_n304), .Y(dp.alu._abc_6356_n458_1) );
	NOR2X1 NOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n305), .Y(dp.alu._abc_6356_n459_1) );
	NAND2X1 NAND2X1_169 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n458_1), .B(dp.alu._abc_6356_n459_1), .Y(dp.alu._abc_6356_n460_1) );
	NAND2X1 NAND2X1_170 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n457_1), .B(dp.alu._abc_6356_n460_1), .Y(aluout_11__RAW) );
	AND2X2 AND2X2_31 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_12_), .B(dp.srcb_12_), .Y(dp.alu._abc_6356_n462_1) );
	AND2X2 AND2X2_32 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n462_1), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n463_1) );
	NOR2X1 NOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_12_), .B(dp.srcb_12_), .Y(dp.alu._abc_6356_n464_1) );
	NOR2X1 NOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n464_1), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n465_1) );
	NOR2X1 NOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n463_1), .B(dp.alu._abc_6356_n465_1), .Y(dp.alu._abc_6356_n466_1) );
	NAND2X1 NAND2X1_171 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n306), .Y(dp.alu._abc_6356_n467_1) );
	NOR2X1 NOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n270), .B(dp.alu._abc_6356_n305), .Y(dp.alu._abc_6356_n468_1) );
	OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n467_1), .B(dp.alu._abc_6356_n468_1), .Y(dp.alu._abc_6356_n469_1) );
	NAND2X1 NAND2X1_172 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n466_1), .B(dp.alu._abc_6356_n469_1), .Y(aluout_12__RAW) );
	AND2X2 AND2X2_33 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_13_), .B(dp.srcb_13_), .Y(dp.alu._abc_6356_n471_1) );
	AND2X2 AND2X2_34 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n471_1), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n472_1) );
	NOR2X1 NOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_13_), .B(dp.srcb_13_), .Y(dp.alu._abc_6356_n473_1) );
	NOR2X1 NOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n473_1), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n474_1) );
	NOR2X1 NOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n472_1), .B(dp.alu._abc_6356_n474_1), .Y(dp.alu._abc_6356_n475_1) );
	NAND2X1 NAND2X1_173 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n306), .B(dp.alu._abc_6356_n308), .Y(dp.alu._abc_6356_n476_1) );
	NOR2X1 NOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n309), .Y(dp.alu._abc_6356_n477_1) );
	NAND2X1 NAND2X1_174 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n476_1), .B(dp.alu._abc_6356_n477_1), .Y(dp.alu._abc_6356_n478_1) );
	NAND2X1 NAND2X1_175 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n475_1), .B(dp.alu._abc_6356_n478_1), .Y(aluout_13__RAW) );
	AND2X2 AND2X2_35 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_14_), .B(dp.srcb_14_), .Y(dp.alu._abc_6356_n480_1) );
	AND2X2 AND2X2_36 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n480_1), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n481_1) );
	NOR2X1 NOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_14_), .B(dp.srcb_14_), .Y(dp.alu._abc_6356_n482_1) );
	NOR2X1 NOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n482_1), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n483_1) );
	NOR2X1 NOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n481_1), .B(dp.alu._abc_6356_n483_1), .Y(dp.alu._abc_6356_n484) );
	NAND2X1 NAND2X1_176 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n310), .Y(dp.alu._abc_6356_n485_1) );
	NOR2X1 NOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n269), .B(dp.alu._abc_6356_n309), .Y(dp.alu._abc_6356_n486_1) );
	OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n485_1), .B(dp.alu._abc_6356_n486_1), .Y(dp.alu._abc_6356_n487) );
	NAND2X1 NAND2X1_177 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n484), .B(dp.alu._abc_6356_n487), .Y(aluout_14__RAW) );
	AND2X2 AND2X2_37 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_15_), .B(dp.srcb_15_), .Y(dp.alu._abc_6356_n489_1) );
	AND2X2 AND2X2_38 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n489_1), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n490) );
	NOR2X1 NOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_15_), .B(dp.srcb_15_), .Y(dp.alu._abc_6356_n491_1) );
	NOR2X1 NOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n491_1), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n492_1) );
	NOR2X1 NOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n490), .B(dp.alu._abc_6356_n492_1), .Y(dp.alu._abc_6356_n493) );
	NAND2X1 NAND2X1_178 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n310), .B(dp.alu._abc_6356_n312), .Y(dp.alu._abc_6356_n494_1) );
	NOR2X1 NOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n313), .Y(dp.alu._abc_6356_n495_1) );
	NAND2X1 NAND2X1_179 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n494_1), .B(dp.alu._abc_6356_n495_1), .Y(dp.alu._abc_6356_n496) );
	NAND2X1 NAND2X1_180 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n493), .B(dp.alu._abc_6356_n496), .Y(aluout_15__RAW) );
	AND2X2 AND2X2_39 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_16_), .B(dp.srcb_16_), .Y(dp.alu._abc_6356_n498_1) );
	AND2X2 AND2X2_40 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n498_1), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n499) );
	NOR2X1 NOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_16_), .B(dp.srcb_16_), .Y(dp.alu._abc_6356_n500_1) );
	NOR2X1 NOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n500_1), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n501_1) );
	NOR2X1 NOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n499), .B(dp.alu._abc_6356_n501_1), .Y(dp.alu._abc_6356_n502) );
	NAND2X1 NAND2X1_181 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n314), .Y(dp.alu._abc_6356_n503_1) );
	NOR2X1 NOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n268), .B(dp.alu._abc_6356_n313), .Y(dp.alu._abc_6356_n504_1) );
	OR2X2 OR2X2_9 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n503_1), .B(dp.alu._abc_6356_n504_1), .Y(dp.alu._abc_6356_n505) );
	NAND2X1 NAND2X1_182 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n502), .B(dp.alu._abc_6356_n505), .Y(aluout_16__RAW) );
	AND2X2 AND2X2_41 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_17_), .B(dp.srcb_17_), .Y(dp.alu._abc_6356_n507_1) );
	AND2X2 AND2X2_42 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n507_1), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n508) );
	NOR2X1 NOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_17_), .B(dp.srcb_17_), .Y(dp.alu._abc_6356_n509_1) );
	NOR2X1 NOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n509_1), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n510_1) );
	NOR2X1 NOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n508), .B(dp.alu._abc_6356_n510_1), .Y(dp.alu._abc_6356_n511) );
	NAND2X1 NAND2X1_183 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n314), .B(dp.alu._abc_6356_n316), .Y(dp.alu._abc_6356_n512_1) );
	NOR2X1 NOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n317), .Y(dp.alu._abc_6356_n513_1) );
	NAND2X1 NAND2X1_184 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n512_1), .B(dp.alu._abc_6356_n513_1), .Y(dp.alu._abc_6356_n514) );
	NAND2X1 NAND2X1_185 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n511), .B(dp.alu._abc_6356_n514), .Y(aluout_17__RAW) );
	AND2X2 AND2X2_43 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_18_), .B(dp.srcb_18_), .Y(dp.alu._abc_6356_n516_1) );
	AND2X2 AND2X2_44 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n516_1), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n517) );
	NOR2X1 NOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_18_), .B(dp.srcb_18_), .Y(dp.alu._abc_6356_n518_1) );
	NOR2X1 NOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n518_1), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n519_1) );
	NOR2X1 NOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n517), .B(dp.alu._abc_6356_n519_1), .Y(dp.alu._abc_6356_n520) );
	NAND2X1 NAND2X1_186 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n318), .Y(dp.alu._abc_6356_n521_1) );
	NOR2X1 NOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n267), .B(dp.alu._abc_6356_n317), .Y(dp.alu._abc_6356_n522_1) );
	OR2X2 OR2X2_10 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n521_1), .B(dp.alu._abc_6356_n522_1), .Y(dp.alu._abc_6356_n523) );
	NAND2X1 NAND2X1_187 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n520), .B(dp.alu._abc_6356_n523), .Y(aluout_18__RAW) );
	AND2X2 AND2X2_45 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_19_), .B(dp.srcb_19_), .Y(dp.alu._abc_6356_n525_1) );
	AND2X2 AND2X2_46 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n525_1), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n526) );
	NOR2X1 NOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_19_), .B(dp.srcb_19_), .Y(dp.alu._abc_6356_n527_1) );
	NOR2X1 NOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n527_1), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n528_1) );
	NOR2X1 NOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n526), .B(dp.alu._abc_6356_n528_1), .Y(dp.alu._abc_6356_n529) );
	NAND2X1 NAND2X1_188 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n318), .B(dp.alu._abc_6356_n320), .Y(dp.alu._abc_6356_n530) );
	NOR2X1 NOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n321), .Y(dp.alu._abc_6356_n531) );
	NAND2X1 NAND2X1_189 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n530), .B(dp.alu._abc_6356_n531), .Y(dp.alu._abc_6356_n532) );
	NAND2X1 NAND2X1_190 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n529), .B(dp.alu._abc_6356_n532), .Y(aluout_19__RAW) );
	AND2X2 AND2X2_47 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_20_), .B(dp.srcb_20_), .Y(dp.alu._abc_6356_n534) );
	AND2X2 AND2X2_48 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n534), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n535) );
	NOR2X1 NOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_20_), .B(dp.srcb_20_), .Y(dp.alu._abc_6356_n536) );
	NOR2X1 NOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n536), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n537) );
	NOR2X1 NOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n535), .B(dp.alu._abc_6356_n537), .Y(dp.alu._abc_6356_n538) );
	NAND2X1 NAND2X1_191 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n322), .Y(dp.alu._abc_6356_n539) );
	NOR2X1 NOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n266), .B(dp.alu._abc_6356_n321), .Y(dp.alu._abc_6356_n540) );
	OR2X2 OR2X2_11 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n539), .B(dp.alu._abc_6356_n540), .Y(dp.alu._abc_6356_n541) );
	NAND2X1 NAND2X1_192 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n538), .B(dp.alu._abc_6356_n541), .Y(aluout_20__RAW) );
	AND2X2 AND2X2_49 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_21_), .B(dp.srcb_21_), .Y(dp.alu._abc_6356_n543) );
	AND2X2 AND2X2_50 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n543), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n544) );
	NOR2X1 NOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_21_), .B(dp.srcb_21_), .Y(dp.alu._abc_6356_n545) );
	NOR2X1 NOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n545), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n546) );
	NOR2X1 NOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n544), .B(dp.alu._abc_6356_n546), .Y(dp.alu._abc_6356_n547) );
	NAND2X1 NAND2X1_193 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n322), .B(dp.alu._abc_6356_n324), .Y(dp.alu._abc_6356_n548) );
	NOR2X1 NOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n325), .Y(dp.alu._abc_6356_n549) );
	NAND2X1 NAND2X1_194 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n548), .B(dp.alu._abc_6356_n549), .Y(dp.alu._abc_6356_n550) );
	NAND2X1 NAND2X1_195 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n547), .B(dp.alu._abc_6356_n550), .Y(aluout_21__RAW) );
	AND2X2 AND2X2_51 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_22_), .B(dp.srcb_22_), .Y(dp.alu._abc_6356_n552) );
	AND2X2 AND2X2_52 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n552), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n553) );
	NOR2X1 NOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_22_), .B(dp.srcb_22_), .Y(dp.alu._abc_6356_n554) );
	NOR2X1 NOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n554), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n555) );
	NOR2X1 NOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n553), .B(dp.alu._abc_6356_n555), .Y(dp.alu._abc_6356_n556) );
	NAND2X1 NAND2X1_196 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n326), .Y(dp.alu._abc_6356_n557) );
	NOR2X1 NOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n265), .B(dp.alu._abc_6356_n325), .Y(dp.alu._abc_6356_n558) );
	OR2X2 OR2X2_12 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n557), .B(dp.alu._abc_6356_n558), .Y(dp.alu._abc_6356_n559) );
	NAND2X1 NAND2X1_197 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n556), .B(dp.alu._abc_6356_n559), .Y(aluout_22__RAW) );
	AND2X2 AND2X2_53 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_23_), .B(dp.srcb_23_), .Y(dp.alu._abc_6356_n561) );
	AND2X2 AND2X2_54 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n561), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n562) );
	NOR2X1 NOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_23_), .B(dp.srcb_23_), .Y(dp.alu._abc_6356_n563) );
	NOR2X1 NOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n563), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n564) );
	NOR2X1 NOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n562), .B(dp.alu._abc_6356_n564), .Y(dp.alu._abc_6356_n565) );
	NAND2X1 NAND2X1_198 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n326), .B(dp.alu._abc_6356_n328), .Y(dp.alu._abc_6356_n566) );
	NOR2X1 NOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n329), .Y(dp.alu._abc_6356_n567) );
	NAND2X1 NAND2X1_199 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n566), .B(dp.alu._abc_6356_n567), .Y(dp.alu._abc_6356_n568) );
	NAND2X1 NAND2X1_200 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n565), .B(dp.alu._abc_6356_n568), .Y(aluout_23__RAW) );
	AND2X2 AND2X2_55 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_24_), .B(dp.srcb_24_), .Y(dp.alu._abc_6356_n570) );
	AND2X2 AND2X2_56 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n570), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n571) );
	NOR2X1 NOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_24_), .B(dp.srcb_24_), .Y(dp.alu._abc_6356_n572) );
	NOR2X1 NOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n572), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n573) );
	NOR2X1 NOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n571), .B(dp.alu._abc_6356_n573), .Y(dp.alu._abc_6356_n574) );
	NAND2X1 NAND2X1_201 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n330), .Y(dp.alu._abc_6356_n575) );
	NOR2X1 NOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n264), .B(dp.alu._abc_6356_n329), .Y(dp.alu._abc_6356_n576) );
	OR2X2 OR2X2_13 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n575), .B(dp.alu._abc_6356_n576), .Y(dp.alu._abc_6356_n577) );
	NAND2X1 NAND2X1_202 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n574), .B(dp.alu._abc_6356_n577), .Y(aluout_24__RAW) );
	AND2X2 AND2X2_57 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_25_), .B(dp.srcb_25_), .Y(dp.alu._abc_6356_n579) );
	AND2X2 AND2X2_58 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n579), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n580) );
	NOR2X1 NOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_25_), .B(dp.srcb_25_), .Y(dp.alu._abc_6356_n581) );
	NOR2X1 NOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n581), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n582) );
	NOR2X1 NOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n580), .B(dp.alu._abc_6356_n582), .Y(dp.alu._abc_6356_n583) );
	NAND2X1 NAND2X1_203 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n330), .B(dp.alu._abc_6356_n332), .Y(dp.alu._abc_6356_n584) );
	NOR2X1 NOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n333), .Y(dp.alu._abc_6356_n585) );
	NAND2X1 NAND2X1_204 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n584), .B(dp.alu._abc_6356_n585), .Y(dp.alu._abc_6356_n586) );
	NAND2X1 NAND2X1_205 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n583), .B(dp.alu._abc_6356_n586), .Y(aluout_25__RAW) );
	AND2X2 AND2X2_59 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_26_), .B(dp.srcb_26_), .Y(dp.alu._abc_6356_n588) );
	AND2X2 AND2X2_60 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n588), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n589) );
	NOR2X1 NOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_26_), .B(dp.srcb_26_), .Y(dp.alu._abc_6356_n590) );
	NOR2X1 NOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n590), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n591) );
	NOR2X1 NOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n589), .B(dp.alu._abc_6356_n591), .Y(dp.alu._abc_6356_n592) );
	NAND2X1 NAND2X1_206 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n334), .Y(dp.alu._abc_6356_n593) );
	NOR2X1 NOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n263), .B(dp.alu._abc_6356_n333), .Y(dp.alu._abc_6356_n594) );
	OR2X2 OR2X2_14 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n593), .B(dp.alu._abc_6356_n594), .Y(dp.alu._abc_6356_n595) );
	NAND2X1 NAND2X1_207 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n592), .B(dp.alu._abc_6356_n595), .Y(aluout_26__RAW) );
	XOR2X1 XOR2X1_84 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n262), .B(dp.alu._abc_6356_n334), .Y(dp.alu._abc_6356_n597) );
	NAND2X1 NAND2X1_208 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n597), .Y(dp.alu._abc_6356_n598) );
	AND2X2 AND2X2_61 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_27_), .B(dp.srcb_27_), .Y(dp.alu._abc_6356_n599) );
	AND2X2 AND2X2_62 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n599), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n600) );
	NOR2X1 NOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_27_), .B(dp.srcb_27_), .Y(dp.alu._abc_6356_n601) );
	NOR2X1 NOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n601), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n602) );
	NOR2X1 NOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n600), .B(dp.alu._abc_6356_n602), .Y(dp.alu._abc_6356_n603) );
	AND2X2 AND2X2_63 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n598), .B(dp.alu._abc_6356_n603), .Y(dp.alu._abc_6356_n604) );
	INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n604), .Y(aluout_27__RAW) );
	AND2X2 AND2X2_64 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_28_), .B(dp.srcb_28_), .Y(dp.alu._abc_6356_n606) );
	AND2X2 AND2X2_65 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n606), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n607) );
	NOR2X1 NOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_28_), .B(dp.srcb_28_), .Y(dp.alu._abc_6356_n608) );
	NOR2X1 NOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n608), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n609) );
	NOR2X1 NOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n607), .B(dp.alu._abc_6356_n609), .Y(dp.alu._abc_6356_n610) );
	XOR2X1 XOR2X1_85 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n261), .B(dp.alu._abc_6356_n335), .Y(dp.alu._abc_6356_n611) );
	NAND2X1 NAND2X1_209 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n611), .Y(dp.alu._abc_6356_n612) );
	NAND2X1 NAND2X1_210 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n610), .B(dp.alu._abc_6356_n612), .Y(aluout_28__RAW) );
	XOR2X1 XOR2X1_86 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n260), .B(dp.alu._abc_6356_n336), .Y(dp.alu._abc_6356_n614_1) );
	NAND2X1 NAND2X1_211 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n614_1), .Y(dp.alu._abc_6356_n615) );
	AND2X2 AND2X2_66 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_29_), .B(dp.srcb_29_), .Y(dp.alu._abc_6356_n616) );
	AND2X2 AND2X2_67 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n616), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n617) );
	NOR2X1 NOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_29_), .B(dp.srcb_29_), .Y(dp.alu._abc_6356_n618) );
	NOR2X1 NOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n618), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n619) );
	NOR2X1 NOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n617), .B(dp.alu._abc_6356_n619), .Y(dp.alu._abc_6356_n620) );
	AND2X2 AND2X2_68 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n615), .B(dp.alu._abc_6356_n620), .Y(dp.alu._abc_6356_n621) );
	INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n621), .Y(aluout_29__RAW) );
	AND2X2 AND2X2_69 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_30_), .B(dp.srcb_30_), .Y(dp.alu._abc_6356_n623) );
	AND2X2 AND2X2_70 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n623), .B(dp.alu._abc_6356_n100), .Y(dp.alu._abc_6356_n624) );
	NOR2X1 NOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(dp.srca_30_), .B(dp.srcb_30_), .Y(dp.alu._abc_6356_n625) );
	NOR2X1 NOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n625), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n626) );
	NOR2X1 NOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n624), .B(dp.alu._abc_6356_n626), .Y(dp.alu._abc_6356_n627) );
	NAND2X1 NAND2X1_212 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n337), .B(dp.alu._abc_6356_n343), .Y(dp.alu._abc_6356_n628) );
	NOR2X1 NOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n104), .B(dp.alu._abc_6356_n344), .Y(dp.alu._abc_6356_n629) );
	NAND2X1 NAND2X1_213 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n628), .B(dp.alu._abc_6356_n629), .Y(dp.alu._abc_6356_n630) );
	NAND2X1 NAND2X1_214 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n627), .B(dp.alu._abc_6356_n630), .Y(aluout_30__RAW) );
	NOR2X1 NOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(alucontrol_1_), .B(dp.alu._abc_6356_n349), .Y(dp.alu._abc_6356_n632) );
	NOR2X1 NOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n348), .B(dp.alu._abc_6356_n102), .Y(dp.alu._abc_6356_n633) );
	NOR2X1 NOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n632), .B(dp.alu._abc_6356_n633), .Y(dp.alu._abc_6356_n634) );
	NAND2X1 NAND2X1_215 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n103_1), .B(dp.alu._abc_6356_n359), .Y(dp.alu._abc_6356_n635) );
	NAND2X1 NAND2X1_216 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n634), .B(dp.alu._abc_6356_n635), .Y(aluout_31__RAW) );
	OR2X2 OR2X2_15 ( .gnd(gnd), .vdd(vdd), .A(aluout[3]), .B(aluout_2__RAW), .Y(dp.alu._abc_6356_n637) );
	OR2X2 OR2X2_16 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n637), .B(aluout_4__RAW), .Y(dp.alu._abc_6356_n638) );
	OR2X2 OR2X2_17 ( .gnd(gnd), .vdd(vdd), .A(aluout_5__RAW), .B(dp.alu._abc_6356_n638), .Y(dp.alu._abc_6356_n639) );
	OR2X2 OR2X2_18 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n639), .B(aluout_6__RAW), .Y(dp.alu._abc_6356_n640) );
	OR2X2 OR2X2_19 ( .gnd(gnd), .vdd(vdd), .A(aluout_7__RAW), .B(dp.alu._abc_6356_n640), .Y(dp.alu._abc_6356_n641) );
	OR2X2 OR2X2_20 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n641), .B(aluout_8__RAW), .Y(dp.alu._abc_6356_n642) );
	OR2X2 OR2X2_21 ( .gnd(gnd), .vdd(vdd), .A(aluout_9__RAW), .B(dp.alu._abc_6356_n642), .Y(dp.alu._abc_6356_n643) );
	NOR2X1 NOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(aluout_10__RAW), .B(dp.alu._abc_6356_n643), .Y(dp.alu._abc_6356_n644) );
	NOR2X1 NOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(aluout_1__RAW), .B(aluout_11__RAW), .Y(dp.alu._abc_6356_n645) );
	NAND2X1 NAND2X1_217 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n644), .B(dp.alu._abc_6356_n645), .Y(dp.alu._abc_6356_n646) );
	OR2X2 OR2X2_22 ( .gnd(gnd), .vdd(vdd), .A(aluout_13__RAW), .B(dp.alu._abc_6356_n646), .Y(dp.alu._abc_6356_n647) );
	OR2X2 OR2X2_23 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n647), .B(aluout_14__RAW), .Y(dp.alu._abc_6356_n648) );
	OR2X2 OR2X2_24 ( .gnd(gnd), .vdd(vdd), .A(aluout_15__RAW), .B(dp.alu._abc_6356_n648), .Y(dp.alu._abc_6356_n649) );
	NOR2X1 NOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(aluout_16__RAW), .B(dp.alu._abc_6356_n649), .Y(dp.alu._abc_6356_n650) );
	NOR2X1 NOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(aluout_12__RAW), .B(aluout_17__RAW), .Y(dp.alu._abc_6356_n651) );
	NAND2X1 NAND2X1_218 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n650), .B(dp.alu._abc_6356_n651), .Y(dp.alu._abc_6356_n652) );
	OR2X2 OR2X2_25 ( .gnd(gnd), .vdd(vdd), .A(aluout_19__RAW), .B(dp.alu._abc_6356_n652), .Y(dp.alu._abc_6356_n653) );
	NOR2X1 NOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(aluout_20__RAW), .B(dp.alu._abc_6356_n653), .Y(dp.alu._abc_6356_n654) );
	NOR2X1 NOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(aluout_18__RAW), .B(aluout_21__RAW), .Y(dp.alu._abc_6356_n655) );
	NAND2X1 NAND2X1_219 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n654), .B(dp.alu._abc_6356_n655), .Y(dp.alu._abc_6356_n656) );
	OR2X2 OR2X2_26 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n656), .B(aluout_22__RAW), .Y(dp.alu._abc_6356_n657) );
	OR2X2 OR2X2_27 ( .gnd(gnd), .vdd(vdd), .A(aluout_23__RAW), .B(dp.alu._abc_6356_n657), .Y(dp.alu._abc_6356_n658) );
	OR2X2 OR2X2_28 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n658), .B(aluout_24__RAW), .Y(dp.alu._abc_6356_n659) );
	OR2X2 OR2X2_29 ( .gnd(gnd), .vdd(vdd), .A(aluout_25__RAW), .B(dp.alu._abc_6356_n659), .Y(dp.alu._abc_6356_n660) );
	NOR2X1 NOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(aluout_26__RAW), .B(dp.alu._abc_6356_n660), .Y(dp.alu._abc_6356_n661) );
	NAND2X1 NAND2X1_220 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n661), .B(dp.alu._abc_6356_n604), .Y(dp.alu._abc_6356_n662) );
	NOR2X1 NOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n662), .B(aluout_28__RAW), .Y(dp.alu._abc_6356_n663) );
	NAND2X1 NAND2X1_221 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n663), .B(dp.alu._abc_6356_n621), .Y(dp.alu._abc_6356_n664) );
	NOR2X1 NOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n664), .B(aluout_30__RAW), .Y(dp.alu._abc_6356_n665) );
	NAND2X1 NAND2X1_222 ( .gnd(gnd), .vdd(vdd), .A(dp.alu._abc_6356_n665), .B(dp.alu._abc_6356_n364), .Y(dp.alu._abc_6356_n666) );
	NOR2X1 NOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(aluout_31__RAW), .B(dp.alu._abc_6356_n666), .Y(zero) );
	NOR2X1 NOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(pc_0__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n96_1) );
	AND2X2 AND2X2_71 ( .gnd(gnd), .vdd(vdd), .A(pc_0__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n97_1) );
	NOR2X1 NOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n96_1), .B(dp.pcadd1._abc_6355_n97_1), .Y(dp.pcplus4_0_) );
	NAND2X1 NAND2X1_223 ( .gnd(gnd), .vdd(vdd), .A(pc_9__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n99) );
	XOR2X1 XOR2X1_87 ( .gnd(gnd), .vdd(vdd), .A(pc_9__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n100) );
	NAND2X1 NAND2X1_224 ( .gnd(gnd), .vdd(vdd), .A(pc_8__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n101_1) );
	XOR2X1 XOR2X1_88 ( .gnd(gnd), .vdd(vdd), .A(pc_8__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n102) );
	NAND2X1 NAND2X1_225 ( .gnd(gnd), .vdd(vdd), .A(pc_7__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n103_1) );
	XOR2X1 XOR2X1_89 ( .gnd(gnd), .vdd(vdd), .A(pc_7__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n104_1) );
	NAND2X1 NAND2X1_226 ( .gnd(gnd), .vdd(vdd), .A(pc_6__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n105) );
	XOR2X1 XOR2X1_90 ( .gnd(gnd), .vdd(vdd), .A(pc_6__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n106) );
	NAND2X1 NAND2X1_227 ( .gnd(gnd), .vdd(vdd), .A(pc_5__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n107) );
	XOR2X1 XOR2X1_91 ( .gnd(gnd), .vdd(vdd), .A(pc_5__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n108_1) );
	NAND2X1 NAND2X1_228 ( .gnd(gnd), .vdd(vdd), .A(pc_4__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n109) );
	XOR2X1 XOR2X1_92 ( .gnd(gnd), .vdd(vdd), .A(pc_4__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n110_1) );
	NAND2X1 NAND2X1_229 ( .gnd(gnd), .vdd(vdd), .A(pc_3__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n111_1) );
	XOR2X1 XOR2X1_93 ( .gnd(gnd), .vdd(vdd), .A(pc_3__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n112) );
	NAND2X1 NAND2X1_230 ( .gnd(gnd), .vdd(vdd), .A(pc_2__RAW), .B(vdd), .Y(dp.pcadd1._abc_6355_n113) );
	XOR2X1 XOR2X1_94 ( .gnd(gnd), .vdd(vdd), .A(pc_2__RAW), .B(vdd), .Y(dp.pcadd1._abc_6355_n114) );
	AND2X2 AND2X2_72 ( .gnd(gnd), .vdd(vdd), .A(pc_1__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n115_1) );
	INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n115_1), .Y(dp.pcadd1._abc_6355_n116) );
	NOR2X1 NOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(pc_1__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n117_1) );
	NOR2X1 NOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n117_1), .B(dp.pcadd1._abc_6355_n115_1), .Y(dp.pcadd1._abc_6355_n118_1) );
	NAND2X1 NAND2X1_231 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n97_1), .B(dp.pcadd1._abc_6355_n118_1), .Y(dp.pcadd1._abc_6355_n119) );
	NAND2X1 NAND2X1_232 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n116), .B(dp.pcadd1._abc_6355_n119), .Y(dp.pcadd1._abc_6355_n120) );
	NAND2X1 NAND2X1_233 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n114), .B(dp.pcadd1._abc_6355_n120), .Y(dp.pcadd1._abc_6355_n121) );
	NAND2X1 NAND2X1_234 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n113), .B(dp.pcadd1._abc_6355_n121), .Y(dp.pcadd1._abc_6355_n122_1) );
	NAND2X1 NAND2X1_235 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n112), .B(dp.pcadd1._abc_6355_n122_1), .Y(dp.pcadd1._abc_6355_n123) );
	NAND2X1 NAND2X1_236 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n111_1), .B(dp.pcadd1._abc_6355_n123), .Y(dp.pcadd1._abc_6355_n124_1) );
	NAND2X1 NAND2X1_237 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n110_1), .B(dp.pcadd1._abc_6355_n124_1), .Y(dp.pcadd1._abc_6355_n125_1) );
	NAND2X1 NAND2X1_238 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n109), .B(dp.pcadd1._abc_6355_n125_1), .Y(dp.pcadd1._abc_6355_n126) );
	NAND2X1 NAND2X1_239 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n108_1), .B(dp.pcadd1._abc_6355_n126), .Y(dp.pcadd1._abc_6355_n127) );
	NAND2X1 NAND2X1_240 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n107), .B(dp.pcadd1._abc_6355_n127), .Y(dp.pcadd1._abc_6355_n128) );
	NAND2X1 NAND2X1_241 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n106), .B(dp.pcadd1._abc_6355_n128), .Y(dp.pcadd1._abc_6355_n129_1) );
	NAND2X1 NAND2X1_242 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n105), .B(dp.pcadd1._abc_6355_n129_1), .Y(dp.pcadd1._abc_6355_n130) );
	NAND2X1 NAND2X1_243 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n104_1), .B(dp.pcadd1._abc_6355_n130), .Y(dp.pcadd1._abc_6355_n131_1) );
	NAND2X1 NAND2X1_244 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n103_1), .B(dp.pcadd1._abc_6355_n131_1), .Y(dp.pcadd1._abc_6355_n132_1) );
	NAND2X1 NAND2X1_245 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n102), .B(dp.pcadd1._abc_6355_n132_1), .Y(dp.pcadd1._abc_6355_n133) );
	NAND2X1 NAND2X1_246 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n101_1), .B(dp.pcadd1._abc_6355_n133), .Y(dp.pcadd1._abc_6355_n134) );
	NAND2X1 NAND2X1_247 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n100), .B(dp.pcadd1._abc_6355_n134), .Y(dp.pcadd1._abc_6355_n135) );
	NAND2X1 NAND2X1_248 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n99), .B(dp.pcadd1._abc_6355_n135), .Y(dp.pcadd1._abc_6355_n136_1) );
	XOR2X1 XOR2X1_95 ( .gnd(gnd), .vdd(vdd), .A(pc_10__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n137) );
	XOR2X1 XOR2X1_96 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n136_1), .B(dp.pcadd1._abc_6355_n137), .Y(dp.pcplus4_10_) );
	NAND2X1 NAND2X1_249 ( .gnd(gnd), .vdd(vdd), .A(pc_10__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n139_1) );
	NAND2X1 NAND2X1_250 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n137), .B(dp.pcadd1._abc_6355_n136_1), .Y(dp.pcadd1._abc_6355_n140) );
	NAND2X1 NAND2X1_251 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n139_1), .B(dp.pcadd1._abc_6355_n140), .Y(dp.pcadd1._abc_6355_n141) );
	XOR2X1 XOR2X1_97 ( .gnd(gnd), .vdd(vdd), .A(pc_11__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n142) );
	XOR2X1 XOR2X1_98 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n141), .B(dp.pcadd1._abc_6355_n142), .Y(dp.pcplus4_11_) );
	NAND2X1 NAND2X1_252 ( .gnd(gnd), .vdd(vdd), .A(pc_11__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n144) );
	NAND2X1 NAND2X1_253 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n142), .B(dp.pcadd1._abc_6355_n141), .Y(dp.pcadd1._abc_6355_n145_1) );
	NAND2X1 NAND2X1_254 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n144), .B(dp.pcadd1._abc_6355_n145_1), .Y(dp.pcadd1._abc_6355_n146_1) );
	XOR2X1 XOR2X1_99 ( .gnd(gnd), .vdd(vdd), .A(pc_12__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n147) );
	XOR2X1 XOR2X1_100 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n146_1), .B(dp.pcadd1._abc_6355_n147), .Y(dp.pcplus4_12_) );
	NAND2X1 NAND2X1_255 ( .gnd(gnd), .vdd(vdd), .A(pc_12__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n149) );
	NAND2X1 NAND2X1_256 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n147), .B(dp.pcadd1._abc_6355_n146_1), .Y(dp.pcadd1._abc_6355_n150_1) );
	NAND2X1 NAND2X1_257 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n149), .B(dp.pcadd1._abc_6355_n150_1), .Y(dp.pcadd1._abc_6355_n151) );
	XOR2X1 XOR2X1_101 ( .gnd(gnd), .vdd(vdd), .A(pc_13__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n152_1) );
	XOR2X1 XOR2X1_102 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n151), .B(dp.pcadd1._abc_6355_n152_1), .Y(dp.pcplus4_13_) );
	NAND2X1 NAND2X1_258 ( .gnd(gnd), .vdd(vdd), .A(pc_13__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n154) );
	NAND2X1 NAND2X1_259 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n152_1), .B(dp.pcadd1._abc_6355_n151), .Y(dp.pcadd1._abc_6355_n155) );
	NAND2X1 NAND2X1_260 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n154), .B(dp.pcadd1._abc_6355_n155), .Y(dp.pcadd1._abc_6355_n156) );
	XOR2X1 XOR2X1_103 ( .gnd(gnd), .vdd(vdd), .A(pc_14__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n157_1) );
	XOR2X1 XOR2X1_104 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n156), .B(dp.pcadd1._abc_6355_n157_1), .Y(dp.pcplus4_14_) );
	NAND2X1 NAND2X1_261 ( .gnd(gnd), .vdd(vdd), .A(pc_14__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n159_1) );
	NAND2X1 NAND2X1_262 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n157_1), .B(dp.pcadd1._abc_6355_n156), .Y(dp.pcadd1._abc_6355_n160_1) );
	NAND2X1 NAND2X1_263 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n159_1), .B(dp.pcadd1._abc_6355_n160_1), .Y(dp.pcadd1._abc_6355_n161) );
	XOR2X1 XOR2X1_105 ( .gnd(gnd), .vdd(vdd), .A(pc_15__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n162) );
	XOR2X1 XOR2X1_106 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n161), .B(dp.pcadd1._abc_6355_n162), .Y(dp.pcplus4_15_) );
	NAND2X1 NAND2X1_264 ( .gnd(gnd), .vdd(vdd), .A(pc_15__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n164_1) );
	NAND2X1 NAND2X1_265 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n162), .B(dp.pcadd1._abc_6355_n161), .Y(dp.pcadd1._abc_6355_n165) );
	NAND2X1 NAND2X1_266 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n164_1), .B(dp.pcadd1._abc_6355_n165), .Y(dp.pcadd1._abc_6355_n166_1) );
	XOR2X1 XOR2X1_107 ( .gnd(gnd), .vdd(vdd), .A(pc_16__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n167_1) );
	XOR2X1 XOR2X1_108 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n166_1), .B(dp.pcadd1._abc_6355_n167_1), .Y(dp.pcplus4_16_) );
	NAND2X1 NAND2X1_267 ( .gnd(gnd), .vdd(vdd), .A(pc_16__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n169_1) );
	NAND2X1 NAND2X1_268 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n167_1), .B(dp.pcadd1._abc_6355_n166_1), .Y(dp.pcadd1._abc_6355_n170_1) );
	NAND2X1 NAND2X1_269 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n169_1), .B(dp.pcadd1._abc_6355_n170_1), .Y(dp.pcadd1._abc_6355_n171_1) );
	XOR2X1 XOR2X1_109 ( .gnd(gnd), .vdd(vdd), .A(pc_17__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n172) );
	XOR2X1 XOR2X1_110 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n171_1), .B(dp.pcadd1._abc_6355_n172), .Y(dp.pcplus4_17_) );
	NAND2X1 NAND2X1_270 ( .gnd(gnd), .vdd(vdd), .A(pc_17__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n174) );
	NAND2X1 NAND2X1_271 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n172), .B(dp.pcadd1._abc_6355_n171_1), .Y(dp.pcadd1._abc_6355_n175_1) );
	NAND2X1 NAND2X1_272 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n174), .B(dp.pcadd1._abc_6355_n175_1), .Y(dp.pcadd1._abc_6355_n176) );
	XOR2X1 XOR2X1_111 ( .gnd(gnd), .vdd(vdd), .A(pc_18__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n177_1) );
	XOR2X1 XOR2X1_112 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n176), .B(dp.pcadd1._abc_6355_n177_1), .Y(dp.pcplus4_18_) );
	NAND2X1 NAND2X1_273 ( .gnd(gnd), .vdd(vdd), .A(pc_18__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n179) );
	NAND2X1 NAND2X1_274 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n177_1), .B(dp.pcadd1._abc_6355_n176), .Y(dp.pcadd1._abc_6355_n180) );
	NAND2X1 NAND2X1_275 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n179), .B(dp.pcadd1._abc_6355_n180), .Y(dp.pcadd1._abc_6355_n181) );
	XOR2X1 XOR2X1_113 ( .gnd(gnd), .vdd(vdd), .A(pc_19__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n182_1) );
	XOR2X1 XOR2X1_114 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n181), .B(dp.pcadd1._abc_6355_n182_1), .Y(dp.pcplus4_19_) );
	XOR2X1 XOR2X1_115 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n118_1), .B(dp.pcadd1._abc_6355_n97_1), .Y(dp.pcplus4_1_) );
	NAND2X1 NAND2X1_276 ( .gnd(gnd), .vdd(vdd), .A(pc_19__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n185_1) );
	NAND2X1 NAND2X1_277 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n182_1), .B(dp.pcadd1._abc_6355_n181), .Y(dp.pcadd1._abc_6355_n186) );
	NAND2X1 NAND2X1_278 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n185_1), .B(dp.pcadd1._abc_6355_n186), .Y(dp.pcadd1._abc_6355_n187) );
	XOR2X1 XOR2X1_116 ( .gnd(gnd), .vdd(vdd), .A(pc_20__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n188) );
	XOR2X1 XOR2X1_117 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n187), .B(dp.pcadd1._abc_6355_n188), .Y(dp.pcplus4_20_) );
	NAND2X1 NAND2X1_279 ( .gnd(gnd), .vdd(vdd), .A(pc_20__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n190) );
	NAND2X1 NAND2X1_280 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n188), .B(dp.pcadd1._abc_6355_n187), .Y(dp.pcadd1._abc_6355_n191_1) );
	NAND2X1 NAND2X1_281 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n190), .B(dp.pcadd1._abc_6355_n191_1), .Y(dp.pcadd1._abc_6355_n192_1) );
	XOR2X1 XOR2X1_118 ( .gnd(gnd), .vdd(vdd), .A(pc_21__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n193) );
	XOR2X1 XOR2X1_119 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n192_1), .B(dp.pcadd1._abc_6355_n193), .Y(dp.pcplus4_21_) );
	NAND2X1 NAND2X1_282 ( .gnd(gnd), .vdd(vdd), .A(pc_21__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n195) );
	NAND2X1 NAND2X1_283 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n193), .B(dp.pcadd1._abc_6355_n192_1), .Y(dp.pcadd1._abc_6355_n196_1) );
	NAND2X1 NAND2X1_284 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n195), .B(dp.pcadd1._abc_6355_n196_1), .Y(dp.pcadd1._abc_6355_n197) );
	XOR2X1 XOR2X1_120 ( .gnd(gnd), .vdd(vdd), .A(pc_22__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n198_1) );
	XOR2X1 XOR2X1_121 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n197), .B(dp.pcadd1._abc_6355_n198_1), .Y(dp.pcplus4_22_) );
	NAND2X1 NAND2X1_285 ( .gnd(gnd), .vdd(vdd), .A(pc_22__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n200) );
	NAND2X1 NAND2X1_286 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n198_1), .B(dp.pcadd1._abc_6355_n197), .Y(dp.pcadd1._abc_6355_n201) );
	NAND2X1 NAND2X1_287 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n200), .B(dp.pcadd1._abc_6355_n201), .Y(dp.pcadd1._abc_6355_n202) );
	XOR2X1 XOR2X1_122 ( .gnd(gnd), .vdd(vdd), .A(pc_23__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n203_1) );
	XOR2X1 XOR2X1_123 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n202), .B(dp.pcadd1._abc_6355_n203_1), .Y(dp.pcplus4_23_) );
	NAND2X1 NAND2X1_288 ( .gnd(gnd), .vdd(vdd), .A(pc_23__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n205_1) );
	NAND2X1 NAND2X1_289 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n203_1), .B(dp.pcadd1._abc_6355_n202), .Y(dp.pcadd1._abc_6355_n206_1) );
	NAND2X1 NAND2X1_290 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n205_1), .B(dp.pcadd1._abc_6355_n206_1), .Y(dp.pcadd1._abc_6355_n207) );
	XOR2X1 XOR2X1_124 ( .gnd(gnd), .vdd(vdd), .A(pc_24__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n208) );
	XOR2X1 XOR2X1_125 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n207), .B(dp.pcadd1._abc_6355_n208), .Y(dp.pcplus4_24_) );
	NAND2X1 NAND2X1_291 ( .gnd(gnd), .vdd(vdd), .A(pc_24__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n210_1) );
	NAND2X1 NAND2X1_292 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n208), .B(dp.pcadd1._abc_6355_n207), .Y(dp.pcadd1._abc_6355_n211) );
	NAND2X1 NAND2X1_293 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n210_1), .B(dp.pcadd1._abc_6355_n211), .Y(dp.pcadd1._abc_6355_n212_1) );
	XOR2X1 XOR2X1_126 ( .gnd(gnd), .vdd(vdd), .A(pc_25__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n213_1) );
	XOR2X1 XOR2X1_127 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n212_1), .B(dp.pcadd1._abc_6355_n213_1), .Y(dp.pcplus4_25_) );
	NAND2X1 NAND2X1_294 ( .gnd(gnd), .vdd(vdd), .A(pc_25__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n215) );
	NAND2X1 NAND2X1_295 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n213_1), .B(dp.pcadd1._abc_6355_n212_1), .Y(dp.pcadd1._abc_6355_n216) );
	NAND2X1 NAND2X1_296 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n215), .B(dp.pcadd1._abc_6355_n216), .Y(dp.pcadd1._abc_6355_n217_1) );
	XOR2X1 XOR2X1_128 ( .gnd(gnd), .vdd(vdd), .A(pc_26__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n218) );
	XOR2X1 XOR2X1_129 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n217_1), .B(dp.pcadd1._abc_6355_n218), .Y(dp.pcplus4_26_) );
	NAND2X1 NAND2X1_297 ( .gnd(gnd), .vdd(vdd), .A(pc_26__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n220) );
	NAND2X1 NAND2X1_298 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n218), .B(dp.pcadd1._abc_6355_n217_1), .Y(dp.pcadd1._abc_6355_n221) );
	NAND2X1 NAND2X1_299 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n220), .B(dp.pcadd1._abc_6355_n221), .Y(dp.pcadd1._abc_6355_n222) );
	XOR2X1 XOR2X1_130 ( .gnd(gnd), .vdd(vdd), .A(pc_27__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n223) );
	XOR2X1 XOR2X1_131 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n222), .B(dp.pcadd1._abc_6355_n223), .Y(dp.pcplus4_27_) );
	NAND2X1 NAND2X1_300 ( .gnd(gnd), .vdd(vdd), .A(pc_27__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n225) );
	NAND2X1 NAND2X1_301 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n223), .B(dp.pcadd1._abc_6355_n222), .Y(dp.pcadd1._abc_6355_n226) );
	NAND2X1 NAND2X1_302 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n225), .B(dp.pcadd1._abc_6355_n226), .Y(dp.pcadd1._abc_6355_n227) );
	XOR2X1 XOR2X1_132 ( .gnd(gnd), .vdd(vdd), .A(pc_28__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n228) );
	XOR2X1 XOR2X1_133 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n227), .B(dp.pcadd1._abc_6355_n228), .Y(dp.pcplus4_28_) );
	NAND2X1 NAND2X1_303 ( .gnd(gnd), .vdd(vdd), .A(pc_28__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n230) );
	NAND2X1 NAND2X1_304 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n228), .B(dp.pcadd1._abc_6355_n227), .Y(dp.pcadd1._abc_6355_n231) );
	NAND2X1 NAND2X1_305 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n230), .B(dp.pcadd1._abc_6355_n231), .Y(dp.pcadd1._abc_6355_n232) );
	XOR2X1 XOR2X1_134 ( .gnd(gnd), .vdd(vdd), .A(pc_29__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n233) );
	XOR2X1 XOR2X1_135 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n232), .B(dp.pcadd1._abc_6355_n233), .Y(dp.pcplus4_29_) );
	XOR2X1 XOR2X1_136 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n120), .B(dp.pcadd1._abc_6355_n114), .Y(dp.pcplus4_2_) );
	NAND2X1 NAND2X1_306 ( .gnd(gnd), .vdd(vdd), .A(pc_29__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n236) );
	NAND2X1 NAND2X1_307 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n233), .B(dp.pcadd1._abc_6355_n232), .Y(dp.pcadd1._abc_6355_n237) );
	NAND2X1 NAND2X1_308 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n236), .B(dp.pcadd1._abc_6355_n237), .Y(dp.pcadd1._abc_6355_n238) );
	XOR2X1 XOR2X1_137 ( .gnd(gnd), .vdd(vdd), .A(pc_30__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n239) );
	XOR2X1 XOR2X1_138 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n238), .B(dp.pcadd1._abc_6355_n239), .Y(dp.pcplus4_30_) );
	NAND2X1 NAND2X1_309 ( .gnd(gnd), .vdd(vdd), .A(pc_30__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n241) );
	NAND2X1 NAND2X1_310 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n239), .B(dp.pcadd1._abc_6355_n238), .Y(dp.pcadd1._abc_6355_n242) );
	NAND2X1 NAND2X1_311 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n241), .B(dp.pcadd1._abc_6355_n242), .Y(dp.pcadd1._abc_6355_n243) );
	XNOR2X1 XNOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(pc_31__RAW), .B(gnd), .Y(dp.pcadd1._abc_6355_n244) );
	XNOR2X1 XNOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n243), .B(dp.pcadd1._abc_6355_n244), .Y(dp.pcplus4_31_) );
	XOR2X1 XOR2X1_139 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n122_1), .B(dp.pcadd1._abc_6355_n112), .Y(dp.pcplus4_3_) );
	XOR2X1 XOR2X1_140 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n124_1), .B(dp.pcadd1._abc_6355_n110_1), .Y(dp.pcplus4_4_) );
	XOR2X1 XOR2X1_141 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n126), .B(dp.pcadd1._abc_6355_n108_1), .Y(dp.pcplus4_5_) );
	XOR2X1 XOR2X1_142 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n128), .B(dp.pcadd1._abc_6355_n106), .Y(dp.pcplus4_6_) );
	XOR2X1 XOR2X1_143 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n130), .B(dp.pcadd1._abc_6355_n104_1), .Y(dp.pcplus4_7_) );
	XOR2X1 XOR2X1_144 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n132_1), .B(dp.pcadd1._abc_6355_n102), .Y(dp.pcplus4_8_) );
	XOR2X1 XOR2X1_145 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd1._abc_6355_n134), .B(dp.pcadd1._abc_6355_n100), .Y(dp.pcplus4_9_) );
	NOR2X1 NOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_0_), .B(gnd), .Y(dp.pcadd2._abc_6355_n96_1) );
	AND2X2 AND2X2_73 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_0_), .B(gnd), .Y(dp.pcadd2._abc_6355_n97_1) );
	NOR2X1 NOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n96_1), .B(dp.pcadd2._abc_6355_n97_1), .Y(dp.pcbranch_0_) );
	NAND2X1 NAND2X1_312 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_9_), .B(instr[7]), .Y(dp.pcadd2._abc_6355_n99) );
	XOR2X1 XOR2X1_146 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_9_), .B(instr[7]), .Y(dp.pcadd2._abc_6355_n100) );
	NAND2X1 NAND2X1_313 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_8_), .B(instr[6]), .Y(dp.pcadd2._abc_6355_n101_1) );
	XOR2X1 XOR2X1_147 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_8_), .B(instr[6]), .Y(dp.pcadd2._abc_6355_n102) );
	NAND2X1 NAND2X1_314 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_7_), .B(instr[5]), .Y(dp.pcadd2._abc_6355_n103_1) );
	XOR2X1 XOR2X1_148 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_7_), .B(instr[5]), .Y(dp.pcadd2._abc_6355_n104_1) );
	NAND2X1 NAND2X1_315 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_6_), .B(instr[4]), .Y(dp.pcadd2._abc_6355_n105) );
	XOR2X1 XOR2X1_149 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_6_), .B(instr[4]), .Y(dp.pcadd2._abc_6355_n106) );
	NAND2X1 NAND2X1_316 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_5_), .B(instr[3]), .Y(dp.pcadd2._abc_6355_n107) );
	XOR2X1 XOR2X1_150 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_5_), .B(instr[3]), .Y(dp.pcadd2._abc_6355_n108_1) );
	NAND2X1 NAND2X1_317 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_4_), .B(instr[2]), .Y(dp.pcadd2._abc_6355_n109) );
	XOR2X1 XOR2X1_151 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_4_), .B(instr[2]), .Y(dp.pcadd2._abc_6355_n110_1) );
	NAND2X1 NAND2X1_318 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_3_), .B(instr[1]), .Y(dp.pcadd2._abc_6355_n111_1) );
	XOR2X1 XOR2X1_152 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_3_), .B(instr[1]), .Y(dp.pcadd2._abc_6355_n112) );
	NAND2X1 NAND2X1_319 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_2_), .B(instr[0]), .Y(dp.pcadd2._abc_6355_n113) );
	XOR2X1 XOR2X1_153 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_2_), .B(instr[0]), .Y(dp.pcadd2._abc_6355_n114) );
	AND2X2 AND2X2_74 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_1_), .B(gnd), .Y(dp.pcadd2._abc_6355_n115_1) );
	INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n115_1), .Y(dp.pcadd2._abc_6355_n116) );
	NOR2X1 NOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_1_), .B(gnd), .Y(dp.pcadd2._abc_6355_n117_1) );
	NOR2X1 NOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n117_1), .B(dp.pcadd2._abc_6355_n115_1), .Y(dp.pcadd2._abc_6355_n118_1) );
	NAND2X1 NAND2X1_320 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n97_1), .B(dp.pcadd2._abc_6355_n118_1), .Y(dp.pcadd2._abc_6355_n119) );
	NAND2X1 NAND2X1_321 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n116), .B(dp.pcadd2._abc_6355_n119), .Y(dp.pcadd2._abc_6355_n120) );
	NAND2X1 NAND2X1_322 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n114), .B(dp.pcadd2._abc_6355_n120), .Y(dp.pcadd2._abc_6355_n121) );
	NAND2X1 NAND2X1_323 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n113), .B(dp.pcadd2._abc_6355_n121), .Y(dp.pcadd2._abc_6355_n122_1) );
	NAND2X1 NAND2X1_324 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n112), .B(dp.pcadd2._abc_6355_n122_1), .Y(dp.pcadd2._abc_6355_n123) );
	NAND2X1 NAND2X1_325 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n111_1), .B(dp.pcadd2._abc_6355_n123), .Y(dp.pcadd2._abc_6355_n124_1) );
	NAND2X1 NAND2X1_326 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n110_1), .B(dp.pcadd2._abc_6355_n124_1), .Y(dp.pcadd2._abc_6355_n125_1) );
	NAND2X1 NAND2X1_327 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n109), .B(dp.pcadd2._abc_6355_n125_1), .Y(dp.pcadd2._abc_6355_n126) );
	NAND2X1 NAND2X1_328 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n108_1), .B(dp.pcadd2._abc_6355_n126), .Y(dp.pcadd2._abc_6355_n127) );
	NAND2X1 NAND2X1_329 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n107), .B(dp.pcadd2._abc_6355_n127), .Y(dp.pcadd2._abc_6355_n128) );
	NAND2X1 NAND2X1_330 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n106), .B(dp.pcadd2._abc_6355_n128), .Y(dp.pcadd2._abc_6355_n129_1) );
	NAND2X1 NAND2X1_331 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n105), .B(dp.pcadd2._abc_6355_n129_1), .Y(dp.pcadd2._abc_6355_n130) );
	NAND2X1 NAND2X1_332 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n104_1), .B(dp.pcadd2._abc_6355_n130), .Y(dp.pcadd2._abc_6355_n131_1) );
	NAND2X1 NAND2X1_333 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n103_1), .B(dp.pcadd2._abc_6355_n131_1), .Y(dp.pcadd2._abc_6355_n132_1) );
	NAND2X1 NAND2X1_334 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n102), .B(dp.pcadd2._abc_6355_n132_1), .Y(dp.pcadd2._abc_6355_n133) );
	NAND2X1 NAND2X1_335 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n101_1), .B(dp.pcadd2._abc_6355_n133), .Y(dp.pcadd2._abc_6355_n134) );
	NAND2X1 NAND2X1_336 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n100), .B(dp.pcadd2._abc_6355_n134), .Y(dp.pcadd2._abc_6355_n135) );
	NAND2X1 NAND2X1_337 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n99), .B(dp.pcadd2._abc_6355_n135), .Y(dp.pcadd2._abc_6355_n136_1) );
	XOR2X1 XOR2X1_154 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_10_), .B(instr[8]), .Y(dp.pcadd2._abc_6355_n137) );
	XOR2X1 XOR2X1_155 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n136_1), .B(dp.pcadd2._abc_6355_n137), .Y(dp.pcbranch_10_) );
	NAND2X1 NAND2X1_338 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_10_), .B(instr[8]), .Y(dp.pcadd2._abc_6355_n139_1) );
	NAND2X1 NAND2X1_339 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n137), .B(dp.pcadd2._abc_6355_n136_1), .Y(dp.pcadd2._abc_6355_n140) );
	NAND2X1 NAND2X1_340 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n139_1), .B(dp.pcadd2._abc_6355_n140), .Y(dp.pcadd2._abc_6355_n141) );
	XOR2X1 XOR2X1_156 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_11_), .B(instr[9]), .Y(dp.pcadd2._abc_6355_n142) );
	XOR2X1 XOR2X1_157 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n141), .B(dp.pcadd2._abc_6355_n142), .Y(dp.pcbranch_11_) );
	NAND2X1 NAND2X1_341 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_11_), .B(instr[9]), .Y(dp.pcadd2._abc_6355_n144) );
	NAND2X1 NAND2X1_342 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n142), .B(dp.pcadd2._abc_6355_n141), .Y(dp.pcadd2._abc_6355_n145_1) );
	NAND2X1 NAND2X1_343 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n144), .B(dp.pcadd2._abc_6355_n145_1), .Y(dp.pcadd2._abc_6355_n146_1) );
	XOR2X1 XOR2X1_158 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_12_), .B(instr[10]), .Y(dp.pcadd2._abc_6355_n147) );
	XOR2X1 XOR2X1_159 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n146_1), .B(dp.pcadd2._abc_6355_n147), .Y(dp.pcbranch_12_) );
	NAND2X1 NAND2X1_344 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_12_), .B(instr[10]), .Y(dp.pcadd2._abc_6355_n149) );
	NAND2X1 NAND2X1_345 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n147), .B(dp.pcadd2._abc_6355_n146_1), .Y(dp.pcadd2._abc_6355_n150_1) );
	NAND2X1 NAND2X1_346 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n149), .B(dp.pcadd2._abc_6355_n150_1), .Y(dp.pcadd2._abc_6355_n151) );
	XOR2X1 XOR2X1_160 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_13_), .B(instr[11]), .Y(dp.pcadd2._abc_6355_n152_1) );
	XOR2X1 XOR2X1_161 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n151), .B(dp.pcadd2._abc_6355_n152_1), .Y(dp.pcbranch_13_) );
	NAND2X1 NAND2X1_347 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_13_), .B(instr[11]), .Y(dp.pcadd2._abc_6355_n154) );
	NAND2X1 NAND2X1_348 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n152_1), .B(dp.pcadd2._abc_6355_n151), .Y(dp.pcadd2._abc_6355_n155) );
	NAND2X1 NAND2X1_349 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n154), .B(dp.pcadd2._abc_6355_n155), .Y(dp.pcadd2._abc_6355_n156) );
	XOR2X1 XOR2X1_162 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_14_), .B(instr[12]), .Y(dp.pcadd2._abc_6355_n157_1) );
	XOR2X1 XOR2X1_163 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n156), .B(dp.pcadd2._abc_6355_n157_1), .Y(dp.pcbranch_14_) );
	NAND2X1 NAND2X1_350 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_14_), .B(instr[12]), .Y(dp.pcadd2._abc_6355_n159_1) );
	NAND2X1 NAND2X1_351 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n157_1), .B(dp.pcadd2._abc_6355_n156), .Y(dp.pcadd2._abc_6355_n160_1) );
	NAND2X1 NAND2X1_352 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n159_1), .B(dp.pcadd2._abc_6355_n160_1), .Y(dp.pcadd2._abc_6355_n161) );
	XOR2X1 XOR2X1_164 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_15_), .B(instr[13]), .Y(dp.pcadd2._abc_6355_n162) );
	XOR2X1 XOR2X1_165 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n161), .B(dp.pcadd2._abc_6355_n162), .Y(dp.pcbranch_15_) );
	NAND2X1 NAND2X1_353 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_15_), .B(instr[13]), .Y(dp.pcadd2._abc_6355_n164_1) );
	NAND2X1 NAND2X1_354 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n162), .B(dp.pcadd2._abc_6355_n161), .Y(dp.pcadd2._abc_6355_n165) );
	NAND2X1 NAND2X1_355 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n164_1), .B(dp.pcadd2._abc_6355_n165), .Y(dp.pcadd2._abc_6355_n166_1) );
	XOR2X1 XOR2X1_166 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_16_), .B(instr[14]), .Y(dp.pcadd2._abc_6355_n167_1) );
	XOR2X1 XOR2X1_167 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n166_1), .B(dp.pcadd2._abc_6355_n167_1), .Y(dp.pcbranch_16_) );
	NAND2X1 NAND2X1_356 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_16_), .B(instr[14]), .Y(dp.pcadd2._abc_6355_n169_1) );
	NAND2X1 NAND2X1_357 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n167_1), .B(dp.pcadd2._abc_6355_n166_1), .Y(dp.pcadd2._abc_6355_n170_1) );
	NAND2X1 NAND2X1_358 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n169_1), .B(dp.pcadd2._abc_6355_n170_1), .Y(dp.pcadd2._abc_6355_n171_1) );
	XOR2X1 XOR2X1_168 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_17_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n172) );
	XOR2X1 XOR2X1_169 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n171_1), .B(dp.pcadd2._abc_6355_n172), .Y(dp.pcbranch_17_) );
	NAND2X1 NAND2X1_359 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_17_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n174) );
	NAND2X1 NAND2X1_360 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n172), .B(dp.pcadd2._abc_6355_n171_1), .Y(dp.pcadd2._abc_6355_n175_1) );
	NAND2X1 NAND2X1_361 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n174), .B(dp.pcadd2._abc_6355_n175_1), .Y(dp.pcadd2._abc_6355_n176) );
	XOR2X1 XOR2X1_170 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_18_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n177_1) );
	XOR2X1 XOR2X1_171 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n176), .B(dp.pcadd2._abc_6355_n177_1), .Y(dp.pcbranch_18_) );
	NAND2X1 NAND2X1_362 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_18_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n179) );
	NAND2X1 NAND2X1_363 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n177_1), .B(dp.pcadd2._abc_6355_n176), .Y(dp.pcadd2._abc_6355_n180) );
	NAND2X1 NAND2X1_364 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n179), .B(dp.pcadd2._abc_6355_n180), .Y(dp.pcadd2._abc_6355_n181) );
	XOR2X1 XOR2X1_172 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_19_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n182_1) );
	XOR2X1 XOR2X1_173 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n181), .B(dp.pcadd2._abc_6355_n182_1), .Y(dp.pcbranch_19_) );
	XOR2X1 XOR2X1_174 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n118_1), .B(dp.pcadd2._abc_6355_n97_1), .Y(dp.pcbranch_1_) );
	NAND2X1 NAND2X1_365 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_19_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n185_1) );
	NAND2X1 NAND2X1_366 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n182_1), .B(dp.pcadd2._abc_6355_n181), .Y(dp.pcadd2._abc_6355_n186) );
	NAND2X1 NAND2X1_367 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n185_1), .B(dp.pcadd2._abc_6355_n186), .Y(dp.pcadd2._abc_6355_n187) );
	XOR2X1 XOR2X1_175 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_20_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n188) );
	XOR2X1 XOR2X1_176 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n187), .B(dp.pcadd2._abc_6355_n188), .Y(dp.pcbranch_20_) );
	NAND2X1 NAND2X1_368 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_20_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n190) );
	NAND2X1 NAND2X1_369 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n188), .B(dp.pcadd2._abc_6355_n187), .Y(dp.pcadd2._abc_6355_n191_1) );
	NAND2X1 NAND2X1_370 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n190), .B(dp.pcadd2._abc_6355_n191_1), .Y(dp.pcadd2._abc_6355_n192_1) );
	XOR2X1 XOR2X1_177 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_21_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n193) );
	XOR2X1 XOR2X1_178 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n192_1), .B(dp.pcadd2._abc_6355_n193), .Y(dp.pcbranch_21_) );
	NAND2X1 NAND2X1_371 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_21_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n195) );
	NAND2X1 NAND2X1_372 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n193), .B(dp.pcadd2._abc_6355_n192_1), .Y(dp.pcadd2._abc_6355_n196_1) );
	NAND2X1 NAND2X1_373 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n195), .B(dp.pcadd2._abc_6355_n196_1), .Y(dp.pcadd2._abc_6355_n197) );
	XOR2X1 XOR2X1_179 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_22_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n198_1) );
	XOR2X1 XOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n197), .B(dp.pcadd2._abc_6355_n198_1), .Y(dp.pcbranch_22_) );
	NAND2X1 NAND2X1_374 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_22_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n200) );
	NAND2X1 NAND2X1_375 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n198_1), .B(dp.pcadd2._abc_6355_n197), .Y(dp.pcadd2._abc_6355_n201) );
	NAND2X1 NAND2X1_376 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n200), .B(dp.pcadd2._abc_6355_n201), .Y(dp.pcadd2._abc_6355_n202) );
	XOR2X1 XOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_23_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n203_1) );
	XOR2X1 XOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n202), .B(dp.pcadd2._abc_6355_n203_1), .Y(dp.pcbranch_23_) );
	NAND2X1 NAND2X1_377 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_23_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n205_1) );
	NAND2X1 NAND2X1_378 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n203_1), .B(dp.pcadd2._abc_6355_n202), .Y(dp.pcadd2._abc_6355_n206_1) );
	NAND2X1 NAND2X1_379 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n205_1), .B(dp.pcadd2._abc_6355_n206_1), .Y(dp.pcadd2._abc_6355_n207) );
	XOR2X1 XOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_24_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n208) );
	XOR2X1 XOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n207), .B(dp.pcadd2._abc_6355_n208), .Y(dp.pcbranch_24_) );
	NAND2X1 NAND2X1_380 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_24_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n210_1) );
	NAND2X1 NAND2X1_381 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n208), .B(dp.pcadd2._abc_6355_n207), .Y(dp.pcadd2._abc_6355_n211) );
	NAND2X1 NAND2X1_382 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n210_1), .B(dp.pcadd2._abc_6355_n211), .Y(dp.pcadd2._abc_6355_n212_1) );
	XOR2X1 XOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_25_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n213_1) );
	XOR2X1 XOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n212_1), .B(dp.pcadd2._abc_6355_n213_1), .Y(dp.pcbranch_25_) );
	NAND2X1 NAND2X1_383 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_25_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n215) );
	NAND2X1 NAND2X1_384 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n213_1), .B(dp.pcadd2._abc_6355_n212_1), .Y(dp.pcadd2._abc_6355_n216) );
	NAND2X1 NAND2X1_385 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n215), .B(dp.pcadd2._abc_6355_n216), .Y(dp.pcadd2._abc_6355_n217_1) );
	XOR2X1 XOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_26_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n218) );
	XOR2X1 XOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n217_1), .B(dp.pcadd2._abc_6355_n218), .Y(dp.pcbranch_26_) );
	NAND2X1 NAND2X1_386 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_26_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n220) );
	NAND2X1 NAND2X1_387 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n218), .B(dp.pcadd2._abc_6355_n217_1), .Y(dp.pcadd2._abc_6355_n221) );
	NAND2X1 NAND2X1_388 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n220), .B(dp.pcadd2._abc_6355_n221), .Y(dp.pcadd2._abc_6355_n222) );
	XOR2X1 XOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_27_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n223) );
	XOR2X1 XOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n222), .B(dp.pcadd2._abc_6355_n223), .Y(dp.pcbranch_27_) );
	NAND2X1 NAND2X1_389 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_27_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n225) );
	NAND2X1 NAND2X1_390 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n223), .B(dp.pcadd2._abc_6355_n222), .Y(dp.pcadd2._abc_6355_n226) );
	NAND2X1 NAND2X1_391 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n225), .B(dp.pcadd2._abc_6355_n226), .Y(dp.pcadd2._abc_6355_n227) );
	XOR2X1 XOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_28_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n228) );
	XOR2X1 XOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n227), .B(dp.pcadd2._abc_6355_n228), .Y(dp.pcbranch_28_) );
	NAND2X1 NAND2X1_392 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_28_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n230) );
	NAND2X1 NAND2X1_393 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n228), .B(dp.pcadd2._abc_6355_n227), .Y(dp.pcadd2._abc_6355_n231) );
	NAND2X1 NAND2X1_394 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n230), .B(dp.pcadd2._abc_6355_n231), .Y(dp.pcadd2._abc_6355_n232) );
	XOR2X1 XOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_29_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n233) );
	XOR2X1 XOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n232), .B(dp.pcadd2._abc_6355_n233), .Y(dp.pcbranch_29_) );
	XOR2X1 XOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n120), .B(dp.pcadd2._abc_6355_n114), .Y(dp.pcbranch_2_) );
	NAND2X1 NAND2X1_395 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_29_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n236) );
	NAND2X1 NAND2X1_396 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n233), .B(dp.pcadd2._abc_6355_n232), .Y(dp.pcadd2._abc_6355_n237) );
	NAND2X1 NAND2X1_397 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n236), .B(dp.pcadd2._abc_6355_n237), .Y(dp.pcadd2._abc_6355_n238) );
	XOR2X1 XOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_30_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n239) );
	XOR2X1 XOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n238), .B(dp.pcadd2._abc_6355_n239), .Y(dp.pcbranch_30_) );
	NAND2X1 NAND2X1_398 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_30_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n241) );
	NAND2X1 NAND2X1_399 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n239), .B(dp.pcadd2._abc_6355_n238), .Y(dp.pcadd2._abc_6355_n242) );
	NAND2X1 NAND2X1_400 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n241), .B(dp.pcadd2._abc_6355_n242), .Y(dp.pcadd2._abc_6355_n243) );
	XNOR2X1 XNOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_31_), .B(instr[15]), .Y(dp.pcadd2._abc_6355_n244) );
	XNOR2X1 XNOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n243), .B(dp.pcadd2._abc_6355_n244), .Y(dp.pcbranch_31_) );
	XOR2X1 XOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n122_1), .B(dp.pcadd2._abc_6355_n112), .Y(dp.pcbranch_3_) );
	XOR2X1 XOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n124_1), .B(dp.pcadd2._abc_6355_n110_1), .Y(dp.pcbranch_4_) );
	XOR2X1 XOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n126), .B(dp.pcadd2._abc_6355_n108_1), .Y(dp.pcbranch_5_) );
	XOR2X1 XOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n128), .B(dp.pcadd2._abc_6355_n106), .Y(dp.pcbranch_6_) );
	XOR2X1 XOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n130), .B(dp.pcadd2._abc_6355_n104_1), .Y(dp.pcbranch_7_) );
	XOR2X1 XOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n132_1), .B(dp.pcadd2._abc_6355_n102), .Y(dp.pcbranch_8_) );
	XOR2X1 XOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(dp.pcadd2._abc_6355_n134), .B(dp.pcadd2._abc_6355_n100), .Y(dp.pcbranch_9_) );
	NAND2X1 NAND2X1_401 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbranch_0_), .B(pcsrc), .Y(dp.pcbrmux._abc_6353_n97) );
	INVX8 INVX8_1 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .Y(dp.pcbrmux._abc_6353_n98) );
	NAND2X1 NAND2X1_402 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_0_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n99) );
	NAND2X1 NAND2X1_403 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n97), .B(dp.pcbrmux._abc_6353_n99), .Y(dp.pcnextbr_0_) );
	NAND2X1 NAND2X1_404 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_1_), .Y(dp.pcbrmux._abc_6353_n101) );
	NAND2X1 NAND2X1_405 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_1_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n102) );
	NAND2X1 NAND2X1_406 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n101), .B(dp.pcbrmux._abc_6353_n102), .Y(dp.pcnextbr_1_) );
	NAND2X1 NAND2X1_407 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_2_), .Y(dp.pcbrmux._abc_6353_n104) );
	NAND2X1 NAND2X1_408 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_2_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n105) );
	NAND2X1 NAND2X1_409 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n104), .B(dp.pcbrmux._abc_6353_n105), .Y(dp.pcnextbr_2_) );
	NAND2X1 NAND2X1_410 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_3_), .Y(dp.pcbrmux._abc_6353_n107) );
	NAND2X1 NAND2X1_411 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_3_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n108) );
	NAND2X1 NAND2X1_412 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n107), .B(dp.pcbrmux._abc_6353_n108), .Y(dp.pcnextbr_3_) );
	NAND2X1 NAND2X1_413 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_4_), .Y(dp.pcbrmux._abc_6353_n110) );
	NAND2X1 NAND2X1_414 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_4_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n111) );
	NAND2X1 NAND2X1_415 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n110), .B(dp.pcbrmux._abc_6353_n111), .Y(dp.pcnextbr_4_) );
	NAND2X1 NAND2X1_416 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_5_), .Y(dp.pcbrmux._abc_6353_n113) );
	NAND2X1 NAND2X1_417 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_5_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n114) );
	NAND2X1 NAND2X1_418 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n113), .B(dp.pcbrmux._abc_6353_n114), .Y(dp.pcnextbr_5_) );
	NAND2X1 NAND2X1_419 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_6_), .Y(dp.pcbrmux._abc_6353_n116) );
	NAND2X1 NAND2X1_420 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_6_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n117) );
	NAND2X1 NAND2X1_421 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n116), .B(dp.pcbrmux._abc_6353_n117), .Y(dp.pcnextbr_6_) );
	NAND2X1 NAND2X1_422 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_7_), .Y(dp.pcbrmux._abc_6353_n119) );
	NAND2X1 NAND2X1_423 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_7_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n120) );
	NAND2X1 NAND2X1_424 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n119), .B(dp.pcbrmux._abc_6353_n120), .Y(dp.pcnextbr_7_) );
	NAND2X1 NAND2X1_425 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_8_), .Y(dp.pcbrmux._abc_6353_n122) );
	NAND2X1 NAND2X1_426 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_8_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n123) );
	NAND2X1 NAND2X1_427 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n122), .B(dp.pcbrmux._abc_6353_n123), .Y(dp.pcnextbr_8_) );
	NAND2X1 NAND2X1_428 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_9_), .Y(dp.pcbrmux._abc_6353_n125) );
	NAND2X1 NAND2X1_429 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_9_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n126) );
	NAND2X1 NAND2X1_430 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n125), .B(dp.pcbrmux._abc_6353_n126), .Y(dp.pcnextbr_9_) );
	NAND2X1 NAND2X1_431 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_10_), .Y(dp.pcbrmux._abc_6353_n128) );
	NAND2X1 NAND2X1_432 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_10_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n129) );
	NAND2X1 NAND2X1_433 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n128), .B(dp.pcbrmux._abc_6353_n129), .Y(dp.pcnextbr_10_) );
	NAND2X1 NAND2X1_434 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_11_), .Y(dp.pcbrmux._abc_6353_n131) );
	NAND2X1 NAND2X1_435 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_11_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n132) );
	NAND2X1 NAND2X1_436 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n131), .B(dp.pcbrmux._abc_6353_n132), .Y(dp.pcnextbr_11_) );
	NAND2X1 NAND2X1_437 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_12_), .Y(dp.pcbrmux._abc_6353_n134) );
	NAND2X1 NAND2X1_438 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_12_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n135) );
	NAND2X1 NAND2X1_439 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n134), .B(dp.pcbrmux._abc_6353_n135), .Y(dp.pcnextbr_12_) );
	NAND2X1 NAND2X1_440 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_13_), .Y(dp.pcbrmux._abc_6353_n137) );
	NAND2X1 NAND2X1_441 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_13_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n138) );
	NAND2X1 NAND2X1_442 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n137), .B(dp.pcbrmux._abc_6353_n138), .Y(dp.pcnextbr_13_) );
	NAND2X1 NAND2X1_443 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_14_), .Y(dp.pcbrmux._abc_6353_n140) );
	NAND2X1 NAND2X1_444 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_14_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n141) );
	NAND2X1 NAND2X1_445 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n140), .B(dp.pcbrmux._abc_6353_n141), .Y(dp.pcnextbr_14_) );
	NAND2X1 NAND2X1_446 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_15_), .Y(dp.pcbrmux._abc_6353_n143) );
	NAND2X1 NAND2X1_447 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_15_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n144) );
	NAND2X1 NAND2X1_448 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n143), .B(dp.pcbrmux._abc_6353_n144), .Y(dp.pcnextbr_15_) );
	NAND2X1 NAND2X1_449 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_16_), .Y(dp.pcbrmux._abc_6353_n146) );
	NAND2X1 NAND2X1_450 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_16_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n147) );
	NAND2X1 NAND2X1_451 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n146), .B(dp.pcbrmux._abc_6353_n147), .Y(dp.pcnextbr_16_) );
	NAND2X1 NAND2X1_452 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_17_), .Y(dp.pcbrmux._abc_6353_n149) );
	NAND2X1 NAND2X1_453 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_17_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n150) );
	NAND2X1 NAND2X1_454 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n149), .B(dp.pcbrmux._abc_6353_n150), .Y(dp.pcnextbr_17_) );
	NAND2X1 NAND2X1_455 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_18_), .Y(dp.pcbrmux._abc_6353_n152) );
	NAND2X1 NAND2X1_456 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_18_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n153) );
	NAND2X1 NAND2X1_457 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n152), .B(dp.pcbrmux._abc_6353_n153), .Y(dp.pcnextbr_18_) );
	NAND2X1 NAND2X1_458 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_19_), .Y(dp.pcbrmux._abc_6353_n155) );
	NAND2X1 NAND2X1_459 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_19_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n156) );
	NAND2X1 NAND2X1_460 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n155), .B(dp.pcbrmux._abc_6353_n156), .Y(dp.pcnextbr_19_) );
	NAND2X1 NAND2X1_461 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_20_), .Y(dp.pcbrmux._abc_6353_n158) );
	NAND2X1 NAND2X1_462 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_20_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n159) );
	NAND2X1 NAND2X1_463 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n158), .B(dp.pcbrmux._abc_6353_n159), .Y(dp.pcnextbr_20_) );
	NAND2X1 NAND2X1_464 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_21_), .Y(dp.pcbrmux._abc_6353_n161) );
	NAND2X1 NAND2X1_465 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_21_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n162) );
	NAND2X1 NAND2X1_466 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n161), .B(dp.pcbrmux._abc_6353_n162), .Y(dp.pcnextbr_21_) );
	NAND2X1 NAND2X1_467 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_22_), .Y(dp.pcbrmux._abc_6353_n164) );
	NAND2X1 NAND2X1_468 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_22_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n165) );
	NAND2X1 NAND2X1_469 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n164), .B(dp.pcbrmux._abc_6353_n165), .Y(dp.pcnextbr_22_) );
	NAND2X1 NAND2X1_470 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_23_), .Y(dp.pcbrmux._abc_6353_n167) );
	NAND2X1 NAND2X1_471 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_23_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n168) );
	NAND2X1 NAND2X1_472 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n167), .B(dp.pcbrmux._abc_6353_n168), .Y(dp.pcnextbr_23_) );
	NAND2X1 NAND2X1_473 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_24_), .Y(dp.pcbrmux._abc_6353_n170) );
	NAND2X1 NAND2X1_474 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_24_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n171) );
	NAND2X1 NAND2X1_475 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n170), .B(dp.pcbrmux._abc_6353_n171), .Y(dp.pcnextbr_24_) );
	NAND2X1 NAND2X1_476 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_25_), .Y(dp.pcbrmux._abc_6353_n173) );
	NAND2X1 NAND2X1_477 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_25_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n174) );
	NAND2X1 NAND2X1_478 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n173), .B(dp.pcbrmux._abc_6353_n174), .Y(dp.pcnextbr_25_) );
	NAND2X1 NAND2X1_479 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_26_), .Y(dp.pcbrmux._abc_6353_n176) );
	NAND2X1 NAND2X1_480 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_26_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n177) );
	NAND2X1 NAND2X1_481 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n176), .B(dp.pcbrmux._abc_6353_n177), .Y(dp.pcnextbr_26_) );
	NAND2X1 NAND2X1_482 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_27_), .Y(dp.pcbrmux._abc_6353_n179) );
	NAND2X1 NAND2X1_483 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_27_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n180) );
	NAND2X1 NAND2X1_484 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n179), .B(dp.pcbrmux._abc_6353_n180), .Y(dp.pcnextbr_27_) );
	NAND2X1 NAND2X1_485 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_28_), .Y(dp.pcbrmux._abc_6353_n182) );
	NAND2X1 NAND2X1_486 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_28_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n183) );
	NAND2X1 NAND2X1_487 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n182), .B(dp.pcbrmux._abc_6353_n183), .Y(dp.pcnextbr_28_) );
	NAND2X1 NAND2X1_488 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_29_), .Y(dp.pcbrmux._abc_6353_n185) );
	NAND2X1 NAND2X1_489 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_29_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n186) );
	NAND2X1 NAND2X1_490 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n185), .B(dp.pcbrmux._abc_6353_n186), .Y(dp.pcnextbr_29_) );
	NAND2X1 NAND2X1_491 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_30_), .Y(dp.pcbrmux._abc_6353_n188) );
	NAND2X1 NAND2X1_492 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_30_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n189) );
	NAND2X1 NAND2X1_493 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n188), .B(dp.pcbrmux._abc_6353_n189), .Y(dp.pcnextbr_30_) );
	NAND2X1 NAND2X1_494 ( .gnd(gnd), .vdd(vdd), .A(pcsrc), .B(dp.pcbranch_31_), .Y(dp.pcbrmux._abc_6353_n191) );
	NAND2X1 NAND2X1_495 ( .gnd(gnd), .vdd(vdd), .A(dp.pcplus4_31_), .B(dp.pcbrmux._abc_6353_n98), .Y(dp.pcbrmux._abc_6353_n192) );
	NAND2X1 NAND2X1_496 ( .gnd(gnd), .vdd(vdd), .A(dp.pcbrmux._abc_6353_n191), .B(dp.pcbrmux._abc_6353_n192), .Y(dp.pcnextbr_31_) );
	NAND2X1 NAND2X1_497 ( .gnd(gnd), .vdd(vdd), .A(gnd), .B(c.md.controls_2_), .Y(dp.pcmux._abc_6353_n97) );
	INVX8 INVX8_2 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .Y(dp.pcmux._abc_6353_n98) );
	NAND2X1 NAND2X1_498 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_0_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n99) );
	NAND2X1 NAND2X1_499 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n97), .B(dp.pcmux._abc_6353_n99), .Y(dp.pcnext_0_) );
	NAND2X1 NAND2X1_500 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(gnd), .Y(dp.pcmux._abc_6353_n101) );
	NAND2X1 NAND2X1_501 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_1_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n102) );
	NAND2X1 NAND2X1_502 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n101), .B(dp.pcmux._abc_6353_n102), .Y(dp.pcnext_1_) );
	NAND2X1 NAND2X1_503 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[0]), .Y(dp.pcmux._abc_6353_n104) );
	NAND2X1 NAND2X1_504 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_2_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n105) );
	NAND2X1 NAND2X1_505 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n104), .B(dp.pcmux._abc_6353_n105), .Y(dp.pcnext_2_) );
	NAND2X1 NAND2X1_506 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[1]), .Y(dp.pcmux._abc_6353_n107) );
	NAND2X1 NAND2X1_507 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_3_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n108) );
	NAND2X1 NAND2X1_508 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n107), .B(dp.pcmux._abc_6353_n108), .Y(dp.pcnext_3_) );
	NAND2X1 NAND2X1_509 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[2]), .Y(dp.pcmux._abc_6353_n110) );
	NAND2X1 NAND2X1_510 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_4_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n111) );
	NAND2X1 NAND2X1_511 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n110), .B(dp.pcmux._abc_6353_n111), .Y(dp.pcnext_4_) );
	NAND2X1 NAND2X1_512 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[3]), .Y(dp.pcmux._abc_6353_n113) );
	NAND2X1 NAND2X1_513 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_5_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n114) );
	NAND2X1 NAND2X1_514 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n113), .B(dp.pcmux._abc_6353_n114), .Y(dp.pcnext_5_) );
	NAND2X1 NAND2X1_515 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[4]), .Y(dp.pcmux._abc_6353_n116) );
	NAND2X1 NAND2X1_516 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_6_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n117) );
	NAND2X1 NAND2X1_517 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n116), .B(dp.pcmux._abc_6353_n117), .Y(dp.pcnext_6_) );
	NAND2X1 NAND2X1_518 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[5]), .Y(dp.pcmux._abc_6353_n119) );
	NAND2X1 NAND2X1_519 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_7_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n120) );
	NAND2X1 NAND2X1_520 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n119), .B(dp.pcmux._abc_6353_n120), .Y(dp.pcnext_7_) );
	NAND2X1 NAND2X1_521 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[6]), .Y(dp.pcmux._abc_6353_n122) );
	NAND2X1 NAND2X1_522 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_8_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n123) );
	NAND2X1 NAND2X1_523 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n122), .B(dp.pcmux._abc_6353_n123), .Y(dp.pcnext_8_) );
	NAND2X1 NAND2X1_524 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[7]), .Y(dp.pcmux._abc_6353_n125) );
	NAND2X1 NAND2X1_525 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_9_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n126) );
	NAND2X1 NAND2X1_526 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n125), .B(dp.pcmux._abc_6353_n126), .Y(dp.pcnext_9_) );
	NAND2X1 NAND2X1_527 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[8]), .Y(dp.pcmux._abc_6353_n128) );
	NAND2X1 NAND2X1_528 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_10_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n129) );
	NAND2X1 NAND2X1_529 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n128), .B(dp.pcmux._abc_6353_n129), .Y(dp.pcnext_10_) );
	NAND2X1 NAND2X1_530 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[9]), .Y(dp.pcmux._abc_6353_n131) );
	NAND2X1 NAND2X1_531 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_11_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n132) );
	NAND2X1 NAND2X1_532 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n131), .B(dp.pcmux._abc_6353_n132), .Y(dp.pcnext_11_) );
	NAND2X1 NAND2X1_533 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[10]), .Y(dp.pcmux._abc_6353_n134) );
	NAND2X1 NAND2X1_534 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_12_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n135) );
	NAND2X1 NAND2X1_535 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n134), .B(dp.pcmux._abc_6353_n135), .Y(dp.pcnext_12_) );
	NAND2X1 NAND2X1_536 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[11]), .Y(dp.pcmux._abc_6353_n137) );
	NAND2X1 NAND2X1_537 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_13_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n138) );
	NAND2X1 NAND2X1_538 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n137), .B(dp.pcmux._abc_6353_n138), .Y(dp.pcnext_13_) );
	NAND2X1 NAND2X1_539 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[12]), .Y(dp.pcmux._abc_6353_n140) );
	NAND2X1 NAND2X1_540 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_14_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n141) );
	NAND2X1 NAND2X1_541 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n140), .B(dp.pcmux._abc_6353_n141), .Y(dp.pcnext_14_) );
	NAND2X1 NAND2X1_542 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[13]), .Y(dp.pcmux._abc_6353_n143) );
	NAND2X1 NAND2X1_543 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_15_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n144) );
	NAND2X1 NAND2X1_544 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n143), .B(dp.pcmux._abc_6353_n144), .Y(dp.pcnext_15_) );
	NAND2X1 NAND2X1_545 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[14]), .Y(dp.pcmux._abc_6353_n146) );
	NAND2X1 NAND2X1_546 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_16_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n147) );
	NAND2X1 NAND2X1_547 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n146), .B(dp.pcmux._abc_6353_n147), .Y(dp.pcnext_16_) );
	NAND2X1 NAND2X1_548 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[15]), .Y(dp.pcmux._abc_6353_n149) );
	NAND2X1 NAND2X1_549 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_17_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n150) );
	NAND2X1 NAND2X1_550 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n149), .B(dp.pcmux._abc_6353_n150), .Y(dp.pcnext_17_) );
	NAND2X1 NAND2X1_551 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[16]), .Y(dp.pcmux._abc_6353_n152) );
	NAND2X1 NAND2X1_552 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_18_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n153) );
	NAND2X1 NAND2X1_553 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n152), .B(dp.pcmux._abc_6353_n153), .Y(dp.pcnext_18_) );
	NAND2X1 NAND2X1_554 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[17]), .Y(dp.pcmux._abc_6353_n155) );
	NAND2X1 NAND2X1_555 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_19_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n156) );
	NAND2X1 NAND2X1_556 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n155), .B(dp.pcmux._abc_6353_n156), .Y(dp.pcnext_19_) );
	NAND2X1 NAND2X1_557 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[18]), .Y(dp.pcmux._abc_6353_n158) );
	NAND2X1 NAND2X1_558 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_20_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n159) );
	NAND2X1 NAND2X1_559 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n158), .B(dp.pcmux._abc_6353_n159), .Y(dp.pcnext_20_) );
	NAND2X1 NAND2X1_560 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[19]), .Y(dp.pcmux._abc_6353_n161) );
	NAND2X1 NAND2X1_561 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_21_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n162) );
	NAND2X1 NAND2X1_562 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n161), .B(dp.pcmux._abc_6353_n162), .Y(dp.pcnext_21_) );
	NAND2X1 NAND2X1_563 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[20]), .Y(dp.pcmux._abc_6353_n164) );
	NAND2X1 NAND2X1_564 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_22_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n165) );
	NAND2X1 NAND2X1_565 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n164), .B(dp.pcmux._abc_6353_n165), .Y(dp.pcnext_22_) );
	NAND2X1 NAND2X1_566 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[21]), .Y(dp.pcmux._abc_6353_n167) );
	NAND2X1 NAND2X1_567 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_23_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n168) );
	NAND2X1 NAND2X1_568 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n167), .B(dp.pcmux._abc_6353_n168), .Y(dp.pcnext_23_) );
	NAND2X1 NAND2X1_569 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[22]), .Y(dp.pcmux._abc_6353_n170) );
	NAND2X1 NAND2X1_570 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_24_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n171) );
	NAND2X1 NAND2X1_571 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n170), .B(dp.pcmux._abc_6353_n171), .Y(dp.pcnext_24_) );
	NAND2X1 NAND2X1_572 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[23]), .Y(dp.pcmux._abc_6353_n173) );
	NAND2X1 NAND2X1_573 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_25_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n174) );
	NAND2X1 NAND2X1_574 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n173), .B(dp.pcmux._abc_6353_n174), .Y(dp.pcnext_25_) );
	NAND2X1 NAND2X1_575 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[24]), .Y(dp.pcmux._abc_6353_n176) );
	NAND2X1 NAND2X1_576 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_26_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n177) );
	NAND2X1 NAND2X1_577 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n176), .B(dp.pcmux._abc_6353_n177), .Y(dp.pcnext_26_) );
	NAND2X1 NAND2X1_578 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(instr[25]), .Y(dp.pcmux._abc_6353_n179) );
	NAND2X1 NAND2X1_579 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_27_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n180) );
	NAND2X1 NAND2X1_580 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n179), .B(dp.pcmux._abc_6353_n180), .Y(dp.pcnext_27_) );
	NAND2X1 NAND2X1_581 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(dp.pcplus4_28_), .Y(dp.pcmux._abc_6353_n182) );
	NAND2X1 NAND2X1_582 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_28_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n183) );
	NAND2X1 NAND2X1_583 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n182), .B(dp.pcmux._abc_6353_n183), .Y(dp.pcnext_28_) );
	NAND2X1 NAND2X1_584 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(dp.pcplus4_29_), .Y(dp.pcmux._abc_6353_n185) );
	NAND2X1 NAND2X1_585 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_29_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n186) );
	NAND2X1 NAND2X1_586 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n185), .B(dp.pcmux._abc_6353_n186), .Y(dp.pcnext_29_) );
	NAND2X1 NAND2X1_587 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(dp.pcplus4_30_), .Y(dp.pcmux._abc_6353_n188) );
	NAND2X1 NAND2X1_588 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_30_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n189) );
	NAND2X1 NAND2X1_589 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n188), .B(dp.pcmux._abc_6353_n189), .Y(dp.pcnext_30_) );
	NAND2X1 NAND2X1_590 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .B(dp.pcplus4_31_), .Y(dp.pcmux._abc_6353_n191) );
	NAND2X1 NAND2X1_591 ( .gnd(gnd), .vdd(vdd), .A(dp.pcnextbr_31_), .B(dp.pcmux._abc_6353_n98), .Y(dp.pcmux._abc_6353_n192) );
	NAND2X1 NAND2X1_592 ( .gnd(gnd), .vdd(vdd), .A(dp.pcmux._abc_6353_n191), .B(dp.pcmux._abc_6353_n192), .Y(dp.pcnext_31_) );
	INVX8 INVX8_3 ( .gnd(gnd), .vdd(vdd), .A(reset), .Y(dp.pcreg._abc_6352_n1) );
	DFFSR DFFSR_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_0_), .Q(pc_0__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_1_), .Q(pc_1__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_2_), .Q(pc_2__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_3_), .Q(pc_3__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_4_), .Q(pc_4__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_5_), .Q(pc_5__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_6_), .Q(pc_6__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_7_), .Q(pc_7__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_8_), .Q(pc_8__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_9_), .Q(pc_9__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_10_), .Q(pc_10__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_11_), .Q(pc_11__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_12_), .Q(pc_12__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_13_), .Q(pc_13__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_14_), .Q(pc_14__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_15_), .Q(pc_15__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_16_), .Q(pc_16__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_17_), .Q(pc_17__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_18_), .Q(pc_18__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_19_), .Q(pc_19__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_20_), .Q(pc_20__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_21_), .Q(pc_21__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_22_), .Q(pc_22__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_23_), .Q(pc_23__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_24_), .Q(pc_24__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_25_), .Q(pc_25__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_26_), .Q(pc_26__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_27_), .Q(pc_27__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_28_), .Q(pc_28__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_29_), .Q(pc_29__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_30_), .Q(pc_30__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	DFFSR DFFSR_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.pcnext_31_), .Q(pc_31__RAW), .R(dp.pcreg._abc_6352_n1), .S(vdd) );
	NAND2X1 NAND2X1_593 ( .gnd(gnd), .vdd(vdd), .A(readdata[0]), .B(c.md.controls_3_), .Y(dp.resmux._abc_6353_n97) );
	INVX8 INVX8_4 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .Y(dp.resmux._abc_6353_n98) );
	NAND2X1 NAND2X1_594 ( .gnd(gnd), .vdd(vdd), .A(aluout_0__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n99) );
	NAND2X1 NAND2X1_595 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n97), .B(dp.resmux._abc_6353_n99), .Y(dp.result_0_) );
	NAND2X1 NAND2X1_596 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[1]), .Y(dp.resmux._abc_6353_n101) );
	NAND2X1 NAND2X1_597 ( .gnd(gnd), .vdd(vdd), .A(aluout_1__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n102) );
	NAND2X1 NAND2X1_598 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n101), .B(dp.resmux._abc_6353_n102), .Y(dp.result_1_) );
	NAND2X1 NAND2X1_599 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[2]), .Y(dp.resmux._abc_6353_n104) );
	NAND2X1 NAND2X1_600 ( .gnd(gnd), .vdd(vdd), .A(aluout_2__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n105) );
	NAND2X1 NAND2X1_601 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n104), .B(dp.resmux._abc_6353_n105), .Y(dp.result_2_) );
	NAND2X1 NAND2X1_602 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[3]), .Y(dp.resmux._abc_6353_n107) );
	NAND2X1 NAND2X1_603 ( .gnd(gnd), .vdd(vdd), .A(aluout_3__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n108) );
	NAND2X1 NAND2X1_604 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n107), .B(dp.resmux._abc_6353_n108), .Y(dp.result_3_) );
	NAND2X1 NAND2X1_605 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[4]), .Y(dp.resmux._abc_6353_n110) );
	NAND2X1 NAND2X1_606 ( .gnd(gnd), .vdd(vdd), .A(aluout_4__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n111) );
	NAND2X1 NAND2X1_607 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n110), .B(dp.resmux._abc_6353_n111), .Y(dp.result_4_) );
	NAND2X1 NAND2X1_608 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[5]), .Y(dp.resmux._abc_6353_n113) );
	NAND2X1 NAND2X1_609 ( .gnd(gnd), .vdd(vdd), .A(aluout_5__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n114) );
	NAND2X1 NAND2X1_610 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n113), .B(dp.resmux._abc_6353_n114), .Y(dp.result_5_) );
	NAND2X1 NAND2X1_611 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[6]), .Y(dp.resmux._abc_6353_n116) );
	NAND2X1 NAND2X1_612 ( .gnd(gnd), .vdd(vdd), .A(aluout_6__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n117) );
	NAND2X1 NAND2X1_613 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n116), .B(dp.resmux._abc_6353_n117), .Y(dp.result_6_) );
	NAND2X1 NAND2X1_614 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[7]), .Y(dp.resmux._abc_6353_n119) );
	NAND2X1 NAND2X1_615 ( .gnd(gnd), .vdd(vdd), .A(aluout_7__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n120) );
	NAND2X1 NAND2X1_616 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n119), .B(dp.resmux._abc_6353_n120), .Y(dp.result_7_) );
	NAND2X1 NAND2X1_617 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[8]), .Y(dp.resmux._abc_6353_n122) );
	NAND2X1 NAND2X1_618 ( .gnd(gnd), .vdd(vdd), .A(aluout_8__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n123) );
	NAND2X1 NAND2X1_619 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n122), .B(dp.resmux._abc_6353_n123), .Y(dp.result_8_) );
	NAND2X1 NAND2X1_620 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[9]), .Y(dp.resmux._abc_6353_n125) );
	NAND2X1 NAND2X1_621 ( .gnd(gnd), .vdd(vdd), .A(aluout_9__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n126) );
	NAND2X1 NAND2X1_622 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n125), .B(dp.resmux._abc_6353_n126), .Y(dp.result_9_) );
	NAND2X1 NAND2X1_623 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[10]), .Y(dp.resmux._abc_6353_n128) );
	NAND2X1 NAND2X1_624 ( .gnd(gnd), .vdd(vdd), .A(aluout_10__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n129) );
	NAND2X1 NAND2X1_625 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n128), .B(dp.resmux._abc_6353_n129), .Y(dp.result_10_) );
	NAND2X1 NAND2X1_626 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[11]), .Y(dp.resmux._abc_6353_n131) );
	NAND2X1 NAND2X1_627 ( .gnd(gnd), .vdd(vdd), .A(aluout_11__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n132) );
	NAND2X1 NAND2X1_628 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n131), .B(dp.resmux._abc_6353_n132), .Y(dp.result_11_) );
	NAND2X1 NAND2X1_629 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[12]), .Y(dp.resmux._abc_6353_n134) );
	NAND2X1 NAND2X1_630 ( .gnd(gnd), .vdd(vdd), .A(aluout_12__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n135) );
	NAND2X1 NAND2X1_631 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n134), .B(dp.resmux._abc_6353_n135), .Y(dp.result_12_) );
	NAND2X1 NAND2X1_632 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[13]), .Y(dp.resmux._abc_6353_n137) );
	NAND2X1 NAND2X1_633 ( .gnd(gnd), .vdd(vdd), .A(aluout_13__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n138) );
	NAND2X1 NAND2X1_634 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n137), .B(dp.resmux._abc_6353_n138), .Y(dp.result_13_) );
	NAND2X1 NAND2X1_635 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[14]), .Y(dp.resmux._abc_6353_n140) );
	NAND2X1 NAND2X1_636 ( .gnd(gnd), .vdd(vdd), .A(aluout_14__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n141) );
	NAND2X1 NAND2X1_637 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n140), .B(dp.resmux._abc_6353_n141), .Y(dp.result_14_) );
	NAND2X1 NAND2X1_638 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[15]), .Y(dp.resmux._abc_6353_n143) );
	NAND2X1 NAND2X1_639 ( .gnd(gnd), .vdd(vdd), .A(aluout_15__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n144) );
	NAND2X1 NAND2X1_640 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n143), .B(dp.resmux._abc_6353_n144), .Y(dp.result_15_) );
	NAND2X1 NAND2X1_641 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[16]), .Y(dp.resmux._abc_6353_n146) );
	NAND2X1 NAND2X1_642 ( .gnd(gnd), .vdd(vdd), .A(aluout_16__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n147) );
	NAND2X1 NAND2X1_643 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n146), .B(dp.resmux._abc_6353_n147), .Y(dp.result_16_) );
	NAND2X1 NAND2X1_644 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[17]), .Y(dp.resmux._abc_6353_n149) );
	NAND2X1 NAND2X1_645 ( .gnd(gnd), .vdd(vdd), .A(aluout_17__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n150) );
	NAND2X1 NAND2X1_646 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n149), .B(dp.resmux._abc_6353_n150), .Y(dp.result_17_) );
	NAND2X1 NAND2X1_647 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[18]), .Y(dp.resmux._abc_6353_n152) );
	NAND2X1 NAND2X1_648 ( .gnd(gnd), .vdd(vdd), .A(aluout_18__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n153) );
	NAND2X1 NAND2X1_649 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n152), .B(dp.resmux._abc_6353_n153), .Y(dp.result_18_) );
	NAND2X1 NAND2X1_650 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[19]), .Y(dp.resmux._abc_6353_n155) );
	NAND2X1 NAND2X1_651 ( .gnd(gnd), .vdd(vdd), .A(aluout_19__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n156) );
	NAND2X1 NAND2X1_652 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n155), .B(dp.resmux._abc_6353_n156), .Y(dp.result_19_) );
	NAND2X1 NAND2X1_653 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[20]), .Y(dp.resmux._abc_6353_n158) );
	NAND2X1 NAND2X1_654 ( .gnd(gnd), .vdd(vdd), .A(aluout_20__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n159) );
	NAND2X1 NAND2X1_655 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n158), .B(dp.resmux._abc_6353_n159), .Y(dp.result_20_) );
	NAND2X1 NAND2X1_656 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[21]), .Y(dp.resmux._abc_6353_n161) );
	NAND2X1 NAND2X1_657 ( .gnd(gnd), .vdd(vdd), .A(aluout_21__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n162) );
	NAND2X1 NAND2X1_658 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n161), .B(dp.resmux._abc_6353_n162), .Y(dp.result_21_) );
	NAND2X1 NAND2X1_659 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[22]), .Y(dp.resmux._abc_6353_n164) );
	NAND2X1 NAND2X1_660 ( .gnd(gnd), .vdd(vdd), .A(aluout_22__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n165) );
	NAND2X1 NAND2X1_661 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n164), .B(dp.resmux._abc_6353_n165), .Y(dp.result_22_) );
	NAND2X1 NAND2X1_662 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[23]), .Y(dp.resmux._abc_6353_n167) );
	NAND2X1 NAND2X1_663 ( .gnd(gnd), .vdd(vdd), .A(aluout_23__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n168) );
	NAND2X1 NAND2X1_664 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n167), .B(dp.resmux._abc_6353_n168), .Y(dp.result_23_) );
	NAND2X1 NAND2X1_665 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[24]), .Y(dp.resmux._abc_6353_n170) );
	NAND2X1 NAND2X1_666 ( .gnd(gnd), .vdd(vdd), .A(aluout_24__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n171) );
	NAND2X1 NAND2X1_667 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n170), .B(dp.resmux._abc_6353_n171), .Y(dp.result_24_) );
	NAND2X1 NAND2X1_668 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[25]), .Y(dp.resmux._abc_6353_n173) );
	NAND2X1 NAND2X1_669 ( .gnd(gnd), .vdd(vdd), .A(aluout_25__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n174) );
	NAND2X1 NAND2X1_670 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n173), .B(dp.resmux._abc_6353_n174), .Y(dp.result_25_) );
	NAND2X1 NAND2X1_671 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[26]), .Y(dp.resmux._abc_6353_n176) );
	NAND2X1 NAND2X1_672 ( .gnd(gnd), .vdd(vdd), .A(aluout_26__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n177) );
	NAND2X1 NAND2X1_673 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n176), .B(dp.resmux._abc_6353_n177), .Y(dp.result_26_) );
	NAND2X1 NAND2X1_674 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[27]), .Y(dp.resmux._abc_6353_n179) );
	NAND2X1 NAND2X1_675 ( .gnd(gnd), .vdd(vdd), .A(aluout_27__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n180) );
	NAND2X1 NAND2X1_676 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n179), .B(dp.resmux._abc_6353_n180), .Y(dp.result_27_) );
	NAND2X1 NAND2X1_677 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[28]), .Y(dp.resmux._abc_6353_n182) );
	NAND2X1 NAND2X1_678 ( .gnd(gnd), .vdd(vdd), .A(aluout_28__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n183) );
	NAND2X1 NAND2X1_679 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n182), .B(dp.resmux._abc_6353_n183), .Y(dp.result_28_) );
	NAND2X1 NAND2X1_680 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[29]), .Y(dp.resmux._abc_6353_n185) );
	NAND2X1 NAND2X1_681 ( .gnd(gnd), .vdd(vdd), .A(aluout_29__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n186) );
	NAND2X1 NAND2X1_682 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n185), .B(dp.resmux._abc_6353_n186), .Y(dp.result_29_) );
	NAND2X1 NAND2X1_683 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[30]), .Y(dp.resmux._abc_6353_n188) );
	NAND2X1 NAND2X1_684 ( .gnd(gnd), .vdd(vdd), .A(aluout_30__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n189) );
	NAND2X1 NAND2X1_685 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n188), .B(dp.resmux._abc_6353_n189), .Y(dp.result_30_) );
	NAND2X1 NAND2X1_686 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .B(readdata[31]), .Y(dp.resmux._abc_6353_n191) );
	NAND2X1 NAND2X1_687 ( .gnd(gnd), .vdd(vdd), .A(aluout_31__RAW), .B(dp.resmux._abc_6353_n98), .Y(dp.resmux._abc_6353_n192) );
	NAND2X1 NAND2X1_688 ( .gnd(gnd), .vdd(vdd), .A(dp.resmux._abc_6353_n191), .B(dp.resmux._abc_6353_n192), .Y(dp.result_31_) );
	INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_8_), .Y(dp.rf._abc_6362_n2160) );
	NOR2X1 NOR2X1_180 ( .gnd(gnd), .vdd(vdd), .A(dp.writereg_4_), .B(dp.rf._abc_6362_n2160), .Y(dp.rf._abc_6362_n2161) );
	INVX4 INVX4_2 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2161), .Y(dp.rf._abc_6362_n2162) );
	INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(dp.writereg_0_), .Y(dp.rf._abc_6362_n2163) );
	NOR2X1 NOR2X1_181 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2163), .B(dp.rf._abc_6362_n2160), .Y(dp.rf._abc_6362_n2164) );
	INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(dp.writereg_1_), .Y(dp.rf._abc_6362_n2165) );
	NOR2X1 NOR2X1_182 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2160), .B(dp.rf._abc_6362_n2165), .Y(dp.rf._abc_6362_n2166) );
	NOR2X1 NOR2X1_183 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2164), .B(dp.rf._abc_6362_n2166), .Y(dp.rf._abc_6362_n2167) );
	INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(dp.writereg_2_), .Y(dp.rf._abc_6362_n2168) );
	NOR2X1 NOR2X1_184 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2160), .B(dp.rf._abc_6362_n2168), .Y(dp.rf._abc_6362_n2169) );
	INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(dp.writereg_3_), .Y(dp.rf._abc_6362_n2170) );
	NOR2X1 NOR2X1_185 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2160), .B(dp.rf._abc_6362_n2170), .Y(dp.rf._abc_6362_n2171) );
	NOR2X1 NOR2X1_186 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2169), .B(dp.rf._abc_6362_n2171), .Y(dp.rf._abc_6362_n2172) );
	NAND2X1 NAND2X1_689 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2167), .B(dp.rf._abc_6362_n2172), .Y(dp.rf._abc_6362_n2173) );
	NOR2X1 NOR2X1_187 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n2173), .Y(dp.rf._abc_6362_n2174) );
	NAND2X1 NAND2X1_690 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2175) );
	INVX8 INVX8_5 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2176) );
	NAND2X1 NAND2X1_691 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<0>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2177) );
	NAND2X1 NAND2X1_692 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2175), .B(dp.rf._abc_6362_n2177), .Y(dp.rf._abc_6362_n3031) );
	NAND2X1 NAND2X1_693 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2179) );
	NAND2X1 NAND2X1_694 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<1>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2180) );
	NAND2X1 NAND2X1_695 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2179), .B(dp.rf._abc_6362_n2180), .Y(dp.rf._abc_6362_n3033) );
	NAND2X1 NAND2X1_696 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2182) );
	NAND2X1 NAND2X1_697 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<2>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2183) );
	NAND2X1 NAND2X1_698 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2182), .B(dp.rf._abc_6362_n2183), .Y(dp.rf._abc_6362_n3035) );
	NAND2X1 NAND2X1_699 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2185) );
	NAND2X1 NAND2X1_700 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<3>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2186) );
	NAND2X1 NAND2X1_701 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2185), .B(dp.rf._abc_6362_n2186), .Y(dp.rf._abc_6362_n3037) );
	NAND2X1 NAND2X1_702 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2188) );
	NAND2X1 NAND2X1_703 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<4>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2189) );
	NAND2X1 NAND2X1_704 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2188), .B(dp.rf._abc_6362_n2189), .Y(dp.rf._abc_6362_n3039) );
	NAND2X1 NAND2X1_705 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2191) );
	NAND2X1 NAND2X1_706 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<5>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2192) );
	NAND2X1 NAND2X1_707 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2191), .B(dp.rf._abc_6362_n2192), .Y(dp.rf._abc_6362_n3041) );
	NAND2X1 NAND2X1_708 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2194) );
	NAND2X1 NAND2X1_709 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<6>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2195) );
	NAND2X1 NAND2X1_710 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2194), .B(dp.rf._abc_6362_n2195), .Y(dp.rf._abc_6362_n3043) );
	NAND2X1 NAND2X1_711 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2197) );
	NAND2X1 NAND2X1_712 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<7>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2198) );
	NAND2X1 NAND2X1_713 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2197), .B(dp.rf._abc_6362_n2198), .Y(dp.rf._abc_6362_n3045) );
	NAND2X1 NAND2X1_714 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2200) );
	NAND2X1 NAND2X1_715 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<8>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2201) );
	NAND2X1 NAND2X1_716 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2200), .B(dp.rf._abc_6362_n2201), .Y(dp.rf._abc_6362_n3047) );
	NAND2X1 NAND2X1_717 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2203) );
	NAND2X1 NAND2X1_718 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<9>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2204) );
	NAND2X1 NAND2X1_719 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2203), .B(dp.rf._abc_6362_n2204), .Y(dp.rf._abc_6362_n3049) );
	NAND2X1 NAND2X1_720 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2206) );
	NAND2X1 NAND2X1_721 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<10>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2207) );
	NAND2X1 NAND2X1_722 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2206), .B(dp.rf._abc_6362_n2207), .Y(dp.rf._abc_6362_n3051) );
	NAND2X1 NAND2X1_723 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2209) );
	NAND2X1 NAND2X1_724 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<11>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2210) );
	NAND2X1 NAND2X1_725 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2209), .B(dp.rf._abc_6362_n2210), .Y(dp.rf._abc_6362_n3053) );
	NAND2X1 NAND2X1_726 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2212) );
	NAND2X1 NAND2X1_727 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<12>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2213) );
	NAND2X1 NAND2X1_728 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2212), .B(dp.rf._abc_6362_n2213), .Y(dp.rf._abc_6362_n3055) );
	NAND2X1 NAND2X1_729 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2215) );
	NAND2X1 NAND2X1_730 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<13>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2216) );
	NAND2X1 NAND2X1_731 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2215), .B(dp.rf._abc_6362_n2216), .Y(dp.rf._abc_6362_n3057) );
	NAND2X1 NAND2X1_732 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2218) );
	NAND2X1 NAND2X1_733 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<14>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2219) );
	NAND2X1 NAND2X1_734 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2218), .B(dp.rf._abc_6362_n2219), .Y(dp.rf._abc_6362_n3059) );
	NAND2X1 NAND2X1_735 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2221) );
	NAND2X1 NAND2X1_736 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<15>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2222) );
	NAND2X1 NAND2X1_737 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2221), .B(dp.rf._abc_6362_n2222), .Y(dp.rf._abc_6362_n3061) );
	NAND2X1 NAND2X1_738 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2224) );
	NAND2X1 NAND2X1_739 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<16>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2225) );
	NAND2X1 NAND2X1_740 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2224), .B(dp.rf._abc_6362_n2225), .Y(dp.rf._abc_6362_n3063) );
	NAND2X1 NAND2X1_741 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2227) );
	NAND2X1 NAND2X1_742 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<17>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2228) );
	NAND2X1 NAND2X1_743 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2227), .B(dp.rf._abc_6362_n2228), .Y(dp.rf._abc_6362_n3065) );
	NAND2X1 NAND2X1_744 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2230) );
	NAND2X1 NAND2X1_745 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<18>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2231) );
	NAND2X1 NAND2X1_746 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2230), .B(dp.rf._abc_6362_n2231), .Y(dp.rf._abc_6362_n3067) );
	NAND2X1 NAND2X1_747 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2233) );
	NAND2X1 NAND2X1_748 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<19>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2234) );
	NAND2X1 NAND2X1_749 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2233), .B(dp.rf._abc_6362_n2234), .Y(dp.rf._abc_6362_n3069) );
	NAND2X1 NAND2X1_750 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2236) );
	NAND2X1 NAND2X1_751 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<20>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2237) );
	NAND2X1 NAND2X1_752 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2236), .B(dp.rf._abc_6362_n2237), .Y(dp.rf._abc_6362_n3071) );
	NAND2X1 NAND2X1_753 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2239) );
	NAND2X1 NAND2X1_754 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<21>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2240) );
	NAND2X1 NAND2X1_755 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2239), .B(dp.rf._abc_6362_n2240), .Y(dp.rf._abc_6362_n3073) );
	NAND2X1 NAND2X1_756 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2242) );
	NAND2X1 NAND2X1_757 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<22>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2243) );
	NAND2X1 NAND2X1_758 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2242), .B(dp.rf._abc_6362_n2243), .Y(dp.rf._abc_6362_n3075) );
	NAND2X1 NAND2X1_759 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2245) );
	NAND2X1 NAND2X1_760 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<23>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2246) );
	NAND2X1 NAND2X1_761 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2245), .B(dp.rf._abc_6362_n2246), .Y(dp.rf._abc_6362_n3077) );
	NAND2X1 NAND2X1_762 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2248) );
	NAND2X1 NAND2X1_763 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<24>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2249) );
	NAND2X1 NAND2X1_764 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2248), .B(dp.rf._abc_6362_n2249), .Y(dp.rf._abc_6362_n3079) );
	NAND2X1 NAND2X1_765 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2251) );
	NAND2X1 NAND2X1_766 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<25>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2252) );
	NAND2X1 NAND2X1_767 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2251), .B(dp.rf._abc_6362_n2252), .Y(dp.rf._abc_6362_n3081) );
	NAND2X1 NAND2X1_768 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2254) );
	NAND2X1 NAND2X1_769 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<26>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2255) );
	NAND2X1 NAND2X1_770 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2254), .B(dp.rf._abc_6362_n2255), .Y(dp.rf._abc_6362_n3083) );
	NAND2X1 NAND2X1_771 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2257) );
	NAND2X1 NAND2X1_772 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<27>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2258) );
	NAND2X1 NAND2X1_773 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2257), .B(dp.rf._abc_6362_n2258), .Y(dp.rf._abc_6362_n3085) );
	NAND2X1 NAND2X1_774 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2260) );
	NAND2X1 NAND2X1_775 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<28>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2261) );
	NAND2X1 NAND2X1_776 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2260), .B(dp.rf._abc_6362_n2261), .Y(dp.rf._abc_6362_n3087) );
	NAND2X1 NAND2X1_777 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2263) );
	NAND2X1 NAND2X1_778 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<29>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2264) );
	NAND2X1 NAND2X1_779 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2263), .B(dp.rf._abc_6362_n2264), .Y(dp.rf._abc_6362_n3089) );
	NAND2X1 NAND2X1_780 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2266) );
	NAND2X1 NAND2X1_781 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<30>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2267) );
	NAND2X1 NAND2X1_782 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2266), .B(dp.rf._abc_6362_n2267), .Y(dp.rf._abc_6362_n3091) );
	NAND2X1 NAND2X1_783 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n2174), .Y(dp.rf._abc_6362_n2269) );
	NAND2X1 NAND2X1_784 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<31>), .B(dp.rf._abc_6362_n2176), .Y(dp.rf._abc_6362_n2270) );
	NAND2X1 NAND2X1_785 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2269), .B(dp.rf._abc_6362_n2270), .Y(dp.rf._abc_6362_n3093) );
	NAND2X1 NAND2X1_786 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2163), .B(dp.rf._abc_6362_n2166), .Y(dp.rf._abc_6362_n2272) );
	INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2272), .Y(dp.rf._abc_6362_n2273) );
	INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2171), .Y(dp.rf._abc_6362_n2274) );
	NOR2X1 NOR2X1_188 ( .gnd(gnd), .vdd(vdd), .A(dp.writereg_2_), .B(dp.rf._abc_6362_n2274), .Y(dp.rf._abc_6362_n2275) );
	NAND2X1 NAND2X1_787 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2273), .B(dp.rf._abc_6362_n2275), .Y(dp.rf._abc_6362_n2276) );
	NOR2X1 NOR2X1_189 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n2276), .Y(dp.rf._abc_6362_n2277) );
	NAND2X1 NAND2X1_788 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2278) );
	INVX8 INVX8_6 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2279) );
	NAND2X1 NAND2X1_789 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<0>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2280) );
	NAND2X1 NAND2X1_790 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2278), .B(dp.rf._abc_6362_n2280), .Y(dp.rf._abc_6362_n3094) );
	NAND2X1 NAND2X1_791 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2282) );
	NAND2X1 NAND2X1_792 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<1>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2283) );
	NAND2X1 NAND2X1_793 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2282), .B(dp.rf._abc_6362_n2283), .Y(dp.rf._abc_6362_n3095) );
	NAND2X1 NAND2X1_794 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2285) );
	NAND2X1 NAND2X1_795 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<2>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2286) );
	NAND2X1 NAND2X1_796 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2285), .B(dp.rf._abc_6362_n2286), .Y(dp.rf._abc_6362_n3096) );
	NAND2X1 NAND2X1_797 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2288) );
	NAND2X1 NAND2X1_798 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<3>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2289) );
	NAND2X1 NAND2X1_799 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2288), .B(dp.rf._abc_6362_n2289), .Y(dp.rf._abc_6362_n3097) );
	NAND2X1 NAND2X1_800 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2291) );
	NAND2X1 NAND2X1_801 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<4>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2292) );
	NAND2X1 NAND2X1_802 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2291), .B(dp.rf._abc_6362_n2292), .Y(dp.rf._abc_6362_n3098) );
	NAND2X1 NAND2X1_803 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2294) );
	NAND2X1 NAND2X1_804 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<5>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2295) );
	NAND2X1 NAND2X1_805 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2294), .B(dp.rf._abc_6362_n2295), .Y(dp.rf._abc_6362_n3099) );
	NAND2X1 NAND2X1_806 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2297) );
	NAND2X1 NAND2X1_807 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<6>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2298) );
	NAND2X1 NAND2X1_808 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2297), .B(dp.rf._abc_6362_n2298), .Y(dp.rf._abc_6362_n3100) );
	NAND2X1 NAND2X1_809 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2300) );
	NAND2X1 NAND2X1_810 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<7>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2301) );
	NAND2X1 NAND2X1_811 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2300), .B(dp.rf._abc_6362_n2301), .Y(dp.rf._abc_6362_n3101) );
	NAND2X1 NAND2X1_812 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2303) );
	NAND2X1 NAND2X1_813 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<8>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2304) );
	NAND2X1 NAND2X1_814 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2303), .B(dp.rf._abc_6362_n2304), .Y(dp.rf._abc_6362_n3102) );
	NAND2X1 NAND2X1_815 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2306) );
	NAND2X1 NAND2X1_816 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<9>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2307) );
	NAND2X1 NAND2X1_817 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2306), .B(dp.rf._abc_6362_n2307), .Y(dp.rf._abc_6362_n3103) );
	NAND2X1 NAND2X1_818 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2309) );
	NAND2X1 NAND2X1_819 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<10>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2310) );
	NAND2X1 NAND2X1_820 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2309), .B(dp.rf._abc_6362_n2310), .Y(dp.rf._abc_6362_n3104) );
	NAND2X1 NAND2X1_821 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2312) );
	NAND2X1 NAND2X1_822 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<11>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2313) );
	NAND2X1 NAND2X1_823 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2312), .B(dp.rf._abc_6362_n2313), .Y(dp.rf._abc_6362_n3105) );
	NAND2X1 NAND2X1_824 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2315) );
	NAND2X1 NAND2X1_825 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<12>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2316) );
	NAND2X1 NAND2X1_826 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2315), .B(dp.rf._abc_6362_n2316), .Y(dp.rf._abc_6362_n3106) );
	NAND2X1 NAND2X1_827 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2318) );
	NAND2X1 NAND2X1_828 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<13>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2319) );
	NAND2X1 NAND2X1_829 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2318), .B(dp.rf._abc_6362_n2319), .Y(dp.rf._abc_6362_n3107) );
	NAND2X1 NAND2X1_830 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2321) );
	NAND2X1 NAND2X1_831 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<14>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2322) );
	NAND2X1 NAND2X1_832 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2321), .B(dp.rf._abc_6362_n2322), .Y(dp.rf._abc_6362_n3108) );
	NAND2X1 NAND2X1_833 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2324) );
	NAND2X1 NAND2X1_834 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<15>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2325) );
	NAND2X1 NAND2X1_835 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2324), .B(dp.rf._abc_6362_n2325), .Y(dp.rf._abc_6362_n3109) );
	NAND2X1 NAND2X1_836 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2327) );
	NAND2X1 NAND2X1_837 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<16>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2328) );
	NAND2X1 NAND2X1_838 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2327), .B(dp.rf._abc_6362_n2328), .Y(dp.rf._abc_6362_n3110) );
	NAND2X1 NAND2X1_839 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2330) );
	NAND2X1 NAND2X1_840 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<17>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2331) );
	NAND2X1 NAND2X1_841 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2330), .B(dp.rf._abc_6362_n2331), .Y(dp.rf._abc_6362_n3111) );
	NAND2X1 NAND2X1_842 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2333) );
	NAND2X1 NAND2X1_843 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<18>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2334) );
	NAND2X1 NAND2X1_844 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2333), .B(dp.rf._abc_6362_n2334), .Y(dp.rf._abc_6362_n3112) );
	NAND2X1 NAND2X1_845 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2336) );
	NAND2X1 NAND2X1_846 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<19>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2337) );
	NAND2X1 NAND2X1_847 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2336), .B(dp.rf._abc_6362_n2337), .Y(dp.rf._abc_6362_n3113) );
	NAND2X1 NAND2X1_848 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2339) );
	NAND2X1 NAND2X1_849 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<20>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2340) );
	NAND2X1 NAND2X1_850 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2339), .B(dp.rf._abc_6362_n2340), .Y(dp.rf._abc_6362_n3114) );
	NAND2X1 NAND2X1_851 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2342) );
	NAND2X1 NAND2X1_852 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<21>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2343) );
	NAND2X1 NAND2X1_853 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2342), .B(dp.rf._abc_6362_n2343), .Y(dp.rf._abc_6362_n3115) );
	NAND2X1 NAND2X1_854 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2345) );
	NAND2X1 NAND2X1_855 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<22>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2346) );
	NAND2X1 NAND2X1_856 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2345), .B(dp.rf._abc_6362_n2346), .Y(dp.rf._abc_6362_n3116) );
	NAND2X1 NAND2X1_857 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2348) );
	NAND2X1 NAND2X1_858 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<23>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2349) );
	NAND2X1 NAND2X1_859 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2348), .B(dp.rf._abc_6362_n2349), .Y(dp.rf._abc_6362_n3117) );
	NAND2X1 NAND2X1_860 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2351) );
	NAND2X1 NAND2X1_861 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<24>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2352) );
	NAND2X1 NAND2X1_862 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2351), .B(dp.rf._abc_6362_n2352), .Y(dp.rf._abc_6362_n3118) );
	NAND2X1 NAND2X1_863 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2354) );
	NAND2X1 NAND2X1_864 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<25>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2355) );
	NAND2X1 NAND2X1_865 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2354), .B(dp.rf._abc_6362_n2355), .Y(dp.rf._abc_6362_n3119) );
	NAND2X1 NAND2X1_866 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2357) );
	NAND2X1 NAND2X1_867 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<26>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2358) );
	NAND2X1 NAND2X1_868 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2357), .B(dp.rf._abc_6362_n2358), .Y(dp.rf._abc_6362_n3120) );
	NAND2X1 NAND2X1_869 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2360) );
	NAND2X1 NAND2X1_870 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<27>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2361) );
	NAND2X1 NAND2X1_871 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2360), .B(dp.rf._abc_6362_n2361), .Y(dp.rf._abc_6362_n3121) );
	NAND2X1 NAND2X1_872 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2363) );
	NAND2X1 NAND2X1_873 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<28>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2364) );
	NAND2X1 NAND2X1_874 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2363), .B(dp.rf._abc_6362_n2364), .Y(dp.rf._abc_6362_n3122) );
	NAND2X1 NAND2X1_875 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2366) );
	NAND2X1 NAND2X1_876 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<29>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2367) );
	NAND2X1 NAND2X1_877 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2366), .B(dp.rf._abc_6362_n2367), .Y(dp.rf._abc_6362_n3123) );
	NAND2X1 NAND2X1_878 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2369) );
	NAND2X1 NAND2X1_879 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<30>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2370) );
	NAND2X1 NAND2X1_880 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2369), .B(dp.rf._abc_6362_n2370), .Y(dp.rf._abc_6362_n3124) );
	NAND2X1 NAND2X1_881 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n2277), .Y(dp.rf._abc_6362_n2372) );
	NAND2X1 NAND2X1_882 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<31>), .B(dp.rf._abc_6362_n2279), .Y(dp.rf._abc_6362_n2373) );
	NAND2X1 NAND2X1_883 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2372), .B(dp.rf._abc_6362_n2373), .Y(dp.rf._abc_6362_n3125) );
	INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2164), .Y(dp.rf._abc_6362_n2375) );
	NOR2X1 NOR2X1_190 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2165), .B(dp.rf._abc_6362_n2375), .Y(dp.rf._abc_6362_n2376) );
	NAND2X1 NAND2X1_884 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2275), .B(dp.rf._abc_6362_n2376), .Y(dp.rf._abc_6362_n2377) );
	NOR2X1 NOR2X1_191 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n2377), .Y(dp.rf._abc_6362_n2378) );
	NAND2X1 NAND2X1_885 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2379) );
	INVX8 INVX8_7 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2380) );
	NAND2X1 NAND2X1_886 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<0>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2381) );
	NAND2X1 NAND2X1_887 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2379), .B(dp.rf._abc_6362_n2381), .Y(dp.rf._abc_6362_n3126) );
	NAND2X1 NAND2X1_888 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2383) );
	NAND2X1 NAND2X1_889 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<1>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2384) );
	NAND2X1 NAND2X1_890 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2383), .B(dp.rf._abc_6362_n2384), .Y(dp.rf._abc_6362_n3127) );
	NAND2X1 NAND2X1_891 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2386) );
	NAND2X1 NAND2X1_892 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<2>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2387) );
	NAND2X1 NAND2X1_893 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2386), .B(dp.rf._abc_6362_n2387), .Y(dp.rf._abc_6362_n3128) );
	NAND2X1 NAND2X1_894 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2389) );
	NAND2X1 NAND2X1_895 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<3>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2390) );
	NAND2X1 NAND2X1_896 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2389), .B(dp.rf._abc_6362_n2390), .Y(dp.rf._abc_6362_n3129) );
	NAND2X1 NAND2X1_897 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2392) );
	NAND2X1 NAND2X1_898 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<4>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2393) );
	NAND2X1 NAND2X1_899 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2392), .B(dp.rf._abc_6362_n2393), .Y(dp.rf._abc_6362_n3130) );
	NAND2X1 NAND2X1_900 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2395) );
	NAND2X1 NAND2X1_901 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<5>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2396) );
	NAND2X1 NAND2X1_902 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2395), .B(dp.rf._abc_6362_n2396), .Y(dp.rf._abc_6362_n3131) );
	NAND2X1 NAND2X1_903 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2398) );
	NAND2X1 NAND2X1_904 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<6>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2399) );
	NAND2X1 NAND2X1_905 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2398), .B(dp.rf._abc_6362_n2399), .Y(dp.rf._abc_6362_n3132) );
	NAND2X1 NAND2X1_906 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2401) );
	NAND2X1 NAND2X1_907 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<7>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2402) );
	NAND2X1 NAND2X1_908 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2401), .B(dp.rf._abc_6362_n2402), .Y(dp.rf._abc_6362_n3133) );
	NAND2X1 NAND2X1_909 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2404) );
	NAND2X1 NAND2X1_910 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<8>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2405) );
	NAND2X1 NAND2X1_911 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2404), .B(dp.rf._abc_6362_n2405), .Y(dp.rf._abc_6362_n3134) );
	NAND2X1 NAND2X1_912 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2407) );
	NAND2X1 NAND2X1_913 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<9>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2408) );
	NAND2X1 NAND2X1_914 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2407), .B(dp.rf._abc_6362_n2408), .Y(dp.rf._abc_6362_n3135) );
	NAND2X1 NAND2X1_915 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2410) );
	NAND2X1 NAND2X1_916 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<10>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2411) );
	NAND2X1 NAND2X1_917 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2410), .B(dp.rf._abc_6362_n2411), .Y(dp.rf._abc_6362_n3136) );
	NAND2X1 NAND2X1_918 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2413) );
	NAND2X1 NAND2X1_919 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<11>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2414) );
	NAND2X1 NAND2X1_920 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2413), .B(dp.rf._abc_6362_n2414), .Y(dp.rf._abc_6362_n3137) );
	NAND2X1 NAND2X1_921 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2416) );
	NAND2X1 NAND2X1_922 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<12>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2417) );
	NAND2X1 NAND2X1_923 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2416), .B(dp.rf._abc_6362_n2417), .Y(dp.rf._abc_6362_n3138) );
	NAND2X1 NAND2X1_924 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2419) );
	NAND2X1 NAND2X1_925 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<13>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2420) );
	NAND2X1 NAND2X1_926 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2419), .B(dp.rf._abc_6362_n2420), .Y(dp.rf._abc_6362_n3139) );
	NAND2X1 NAND2X1_927 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2422) );
	NAND2X1 NAND2X1_928 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<14>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2423) );
	NAND2X1 NAND2X1_929 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2422), .B(dp.rf._abc_6362_n2423), .Y(dp.rf._abc_6362_n3140) );
	NAND2X1 NAND2X1_930 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2425) );
	NAND2X1 NAND2X1_931 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<15>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2426) );
	NAND2X1 NAND2X1_932 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2425), .B(dp.rf._abc_6362_n2426), .Y(dp.rf._abc_6362_n3141) );
	NAND2X1 NAND2X1_933 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2428) );
	NAND2X1 NAND2X1_934 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<16>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2429) );
	NAND2X1 NAND2X1_935 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2428), .B(dp.rf._abc_6362_n2429), .Y(dp.rf._abc_6362_n3142) );
	NAND2X1 NAND2X1_936 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2431) );
	NAND2X1 NAND2X1_937 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<17>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2432) );
	NAND2X1 NAND2X1_938 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2431), .B(dp.rf._abc_6362_n2432), .Y(dp.rf._abc_6362_n3143) );
	NAND2X1 NAND2X1_939 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2434) );
	NAND2X1 NAND2X1_940 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<18>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2435) );
	NAND2X1 NAND2X1_941 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2434), .B(dp.rf._abc_6362_n2435), .Y(dp.rf._abc_6362_n3144) );
	NAND2X1 NAND2X1_942 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2437) );
	NAND2X1 NAND2X1_943 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<19>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2438) );
	NAND2X1 NAND2X1_944 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2437), .B(dp.rf._abc_6362_n2438), .Y(dp.rf._abc_6362_n3145) );
	NAND2X1 NAND2X1_945 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2440) );
	NAND2X1 NAND2X1_946 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<20>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2441) );
	NAND2X1 NAND2X1_947 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2440), .B(dp.rf._abc_6362_n2441), .Y(dp.rf._abc_6362_n3146) );
	NAND2X1 NAND2X1_948 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2443) );
	NAND2X1 NAND2X1_949 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<21>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2444) );
	NAND2X1 NAND2X1_950 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2443), .B(dp.rf._abc_6362_n2444), .Y(dp.rf._abc_6362_n3147) );
	NAND2X1 NAND2X1_951 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2446) );
	NAND2X1 NAND2X1_952 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<22>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2447) );
	NAND2X1 NAND2X1_953 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2446), .B(dp.rf._abc_6362_n2447), .Y(dp.rf._abc_6362_n3148) );
	NAND2X1 NAND2X1_954 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2449) );
	NAND2X1 NAND2X1_955 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<23>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2450) );
	NAND2X1 NAND2X1_956 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2449), .B(dp.rf._abc_6362_n2450), .Y(dp.rf._abc_6362_n3149) );
	NAND2X1 NAND2X1_957 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2452) );
	NAND2X1 NAND2X1_958 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<24>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2453) );
	NAND2X1 NAND2X1_959 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2452), .B(dp.rf._abc_6362_n2453), .Y(dp.rf._abc_6362_n3150) );
	NAND2X1 NAND2X1_960 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2455) );
	NAND2X1 NAND2X1_961 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<25>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2456) );
	NAND2X1 NAND2X1_962 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2455), .B(dp.rf._abc_6362_n2456), .Y(dp.rf._abc_6362_n3151) );
	NAND2X1 NAND2X1_963 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2458) );
	NAND2X1 NAND2X1_964 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<26>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2459) );
	NAND2X1 NAND2X1_965 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2458), .B(dp.rf._abc_6362_n2459), .Y(dp.rf._abc_6362_n3152) );
	NAND2X1 NAND2X1_966 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2461) );
	NAND2X1 NAND2X1_967 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<27>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2462) );
	NAND2X1 NAND2X1_968 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2461), .B(dp.rf._abc_6362_n2462), .Y(dp.rf._abc_6362_n3153) );
	NAND2X1 NAND2X1_969 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2464) );
	NAND2X1 NAND2X1_970 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<28>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2465) );
	NAND2X1 NAND2X1_971 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2464), .B(dp.rf._abc_6362_n2465), .Y(dp.rf._abc_6362_n3154) );
	NAND2X1 NAND2X1_972 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2467) );
	NAND2X1 NAND2X1_973 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<29>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2468) );
	NAND2X1 NAND2X1_974 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2467), .B(dp.rf._abc_6362_n2468), .Y(dp.rf._abc_6362_n3155) );
	NAND2X1 NAND2X1_975 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2470) );
	NAND2X1 NAND2X1_976 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<30>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2471) );
	NAND2X1 NAND2X1_977 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2470), .B(dp.rf._abc_6362_n2471), .Y(dp.rf._abc_6362_n3156) );
	NAND2X1 NAND2X1_978 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n2378), .Y(dp.rf._abc_6362_n2473) );
	NAND2X1 NAND2X1_979 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_11_<31>), .B(dp.rf._abc_6362_n2380), .Y(dp.rf._abc_6362_n2474) );
	NAND2X1 NAND2X1_980 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2473), .B(dp.rf._abc_6362_n2474), .Y(dp.rf._abc_6362_n3157) );
	NOR2X1 NOR2X1_192 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2168), .B(dp.rf._abc_6362_n2274), .Y(dp.rf._abc_6362_n2476) );
	NAND2X1 NAND2X1_981 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2167), .B(dp.rf._abc_6362_n2476), .Y(dp.rf._abc_6362_n2477) );
	NOR2X1 NOR2X1_193 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n2477), .Y(dp.rf._abc_6362_n2478) );
	NAND2X1 NAND2X1_982 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2479) );
	INVX8 INVX8_8 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2480) );
	NAND2X1 NAND2X1_983 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<0>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2481) );
	NAND2X1 NAND2X1_984 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2479), .B(dp.rf._abc_6362_n2481), .Y(dp.rf._abc_6362_n3158) );
	NAND2X1 NAND2X1_985 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2483) );
	NAND2X1 NAND2X1_986 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<1>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2484) );
	NAND2X1 NAND2X1_987 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2483), .B(dp.rf._abc_6362_n2484), .Y(dp.rf._abc_6362_n3159) );
	NAND2X1 NAND2X1_988 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2486) );
	NAND2X1 NAND2X1_989 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<2>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2487) );
	NAND2X1 NAND2X1_990 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2486), .B(dp.rf._abc_6362_n2487), .Y(dp.rf._abc_6362_n3160) );
	NAND2X1 NAND2X1_991 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2489) );
	NAND2X1 NAND2X1_992 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<3>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2490) );
	NAND2X1 NAND2X1_993 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2489), .B(dp.rf._abc_6362_n2490), .Y(dp.rf._abc_6362_n3161) );
	NAND2X1 NAND2X1_994 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2492) );
	NAND2X1 NAND2X1_995 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<4>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2493) );
	NAND2X1 NAND2X1_996 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2492), .B(dp.rf._abc_6362_n2493), .Y(dp.rf._abc_6362_n3162) );
	NAND2X1 NAND2X1_997 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2495) );
	NAND2X1 NAND2X1_998 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<5>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2496) );
	NAND2X1 NAND2X1_999 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2495), .B(dp.rf._abc_6362_n2496), .Y(dp.rf._abc_6362_n3163) );
	NAND2X1 NAND2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2498) );
	NAND2X1 NAND2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<6>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2499) );
	NAND2X1 NAND2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2498), .B(dp.rf._abc_6362_n2499), .Y(dp.rf._abc_6362_n3164) );
	NAND2X1 NAND2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2501) );
	NAND2X1 NAND2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<7>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2502) );
	NAND2X1 NAND2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2501), .B(dp.rf._abc_6362_n2502), .Y(dp.rf._abc_6362_n3165) );
	NAND2X1 NAND2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2504) );
	NAND2X1 NAND2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<8>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2505) );
	NAND2X1 NAND2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2504), .B(dp.rf._abc_6362_n2505), .Y(dp.rf._abc_6362_n3166) );
	NAND2X1 NAND2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2507) );
	NAND2X1 NAND2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<9>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2508) );
	NAND2X1 NAND2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2507), .B(dp.rf._abc_6362_n2508), .Y(dp.rf._abc_6362_n3167) );
	NAND2X1 NAND2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2510) );
	NAND2X1 NAND2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<10>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2511) );
	NAND2X1 NAND2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2510), .B(dp.rf._abc_6362_n2511), .Y(dp.rf._abc_6362_n3168) );
	NAND2X1 NAND2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2513) );
	NAND2X1 NAND2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<11>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2514) );
	NAND2X1 NAND2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2513), .B(dp.rf._abc_6362_n2514), .Y(dp.rf._abc_6362_n3169) );
	NAND2X1 NAND2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2516) );
	NAND2X1 NAND2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<12>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2517) );
	NAND2X1 NAND2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2516), .B(dp.rf._abc_6362_n2517), .Y(dp.rf._abc_6362_n3170) );
	NAND2X1 NAND2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2519) );
	NAND2X1 NAND2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<13>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2520) );
	NAND2X1 NAND2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2519), .B(dp.rf._abc_6362_n2520), .Y(dp.rf._abc_6362_n3171) );
	NAND2X1 NAND2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2522) );
	NAND2X1 NAND2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<14>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2523) );
	NAND2X1 NAND2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2522), .B(dp.rf._abc_6362_n2523), .Y(dp.rf._abc_6362_n3172) );
	NAND2X1 NAND2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2525) );
	NAND2X1 NAND2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<15>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2526) );
	NAND2X1 NAND2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2525), .B(dp.rf._abc_6362_n2526), .Y(dp.rf._abc_6362_n3173) );
	NAND2X1 NAND2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2528) );
	NAND2X1 NAND2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<16>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2529) );
	NAND2X1 NAND2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2528), .B(dp.rf._abc_6362_n2529), .Y(dp.rf._abc_6362_n3174) );
	NAND2X1 NAND2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2531) );
	NAND2X1 NAND2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<17>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2532) );
	NAND2X1 NAND2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2531), .B(dp.rf._abc_6362_n2532), .Y(dp.rf._abc_6362_n3175) );
	NAND2X1 NAND2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2534) );
	NAND2X1 NAND2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<18>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2535) );
	NAND2X1 NAND2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2534), .B(dp.rf._abc_6362_n2535), .Y(dp.rf._abc_6362_n3176) );
	NAND2X1 NAND2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2537) );
	NAND2X1 NAND2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<19>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2538) );
	NAND2X1 NAND2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2537), .B(dp.rf._abc_6362_n2538), .Y(dp.rf._abc_6362_n3177) );
	NAND2X1 NAND2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2540) );
	NAND2X1 NAND2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<20>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2541) );
	NAND2X1 NAND2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2540), .B(dp.rf._abc_6362_n2541), .Y(dp.rf._abc_6362_n3178) );
	NAND2X1 NAND2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2543) );
	NAND2X1 NAND2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<21>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2544) );
	NAND2X1 NAND2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2543), .B(dp.rf._abc_6362_n2544), .Y(dp.rf._abc_6362_n3179) );
	NAND2X1 NAND2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2546) );
	NAND2X1 NAND2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<22>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2547) );
	NAND2X1 NAND2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2546), .B(dp.rf._abc_6362_n2547), .Y(dp.rf._abc_6362_n3180) );
	NAND2X1 NAND2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2549) );
	NAND2X1 NAND2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<23>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2550) );
	NAND2X1 NAND2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2549), .B(dp.rf._abc_6362_n2550), .Y(dp.rf._abc_6362_n3181) );
	NAND2X1 NAND2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2552) );
	NAND2X1 NAND2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<24>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2553) );
	NAND2X1 NAND2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2552), .B(dp.rf._abc_6362_n2553), .Y(dp.rf._abc_6362_n3182) );
	NAND2X1 NAND2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2555) );
	NAND2X1 NAND2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<25>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2556) );
	NAND2X1 NAND2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2555), .B(dp.rf._abc_6362_n2556), .Y(dp.rf._abc_6362_n3183) );
	NAND2X1 NAND2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2558) );
	NAND2X1 NAND2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<26>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2559) );
	NAND2X1 NAND2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2558), .B(dp.rf._abc_6362_n2559), .Y(dp.rf._abc_6362_n3184) );
	NAND2X1 NAND2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2561) );
	NAND2X1 NAND2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<27>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2562) );
	NAND2X1 NAND2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2561), .B(dp.rf._abc_6362_n2562), .Y(dp.rf._abc_6362_n3185) );
	NAND2X1 NAND2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2564) );
	NAND2X1 NAND2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<28>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2565) );
	NAND2X1 NAND2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2564), .B(dp.rf._abc_6362_n2565), .Y(dp.rf._abc_6362_n3186) );
	NAND2X1 NAND2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2567) );
	NAND2X1 NAND2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<29>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2568) );
	NAND2X1 NAND2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2567), .B(dp.rf._abc_6362_n2568), .Y(dp.rf._abc_6362_n3187) );
	NAND2X1 NAND2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2570) );
	NAND2X1 NAND2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<30>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2571) );
	NAND2X1 NAND2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2570), .B(dp.rf._abc_6362_n2571), .Y(dp.rf._abc_6362_n3188) );
	NAND2X1 NAND2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n2478), .Y(dp.rf._abc_6362_n2573) );
	NAND2X1 NAND2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<31>), .B(dp.rf._abc_6362_n2480), .Y(dp.rf._abc_6362_n2574) );
	NAND2X1 NAND2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2573), .B(dp.rf._abc_6362_n2574), .Y(dp.rf._abc_6362_n3189) );
	NOR2X1 NOR2X1_194 ( .gnd(gnd), .vdd(vdd), .A(dp.writereg_1_), .B(dp.rf._abc_6362_n2375), .Y(dp.rf._abc_6362_n2576) );
	NAND2X1 NAND2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2476), .B(dp.rf._abc_6362_n2576), .Y(dp.rf._abc_6362_n2577) );
	NOR2X1 NOR2X1_195 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n2577), .Y(dp.rf._abc_6362_n2578) );
	NAND2X1 NAND2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2579) );
	INVX8 INVX8_9 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2580) );
	NAND2X1 NAND2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<0>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2581) );
	NAND2X1 NAND2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2579), .B(dp.rf._abc_6362_n2581), .Y(dp.rf._abc_6362_n3190) );
	NAND2X1 NAND2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2583) );
	NAND2X1 NAND2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<1>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2584) );
	NAND2X1 NAND2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2583), .B(dp.rf._abc_6362_n2584), .Y(dp.rf._abc_6362_n3191) );
	NAND2X1 NAND2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2586) );
	NAND2X1 NAND2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<2>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2587) );
	NAND2X1 NAND2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2586), .B(dp.rf._abc_6362_n2587), .Y(dp.rf._abc_6362_n3192) );
	NAND2X1 NAND2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2589) );
	NAND2X1 NAND2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<3>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2590) );
	NAND2X1 NAND2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2589), .B(dp.rf._abc_6362_n2590), .Y(dp.rf._abc_6362_n3193) );
	NAND2X1 NAND2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2592) );
	NAND2X1 NAND2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<4>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2593) );
	NAND2X1 NAND2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2592), .B(dp.rf._abc_6362_n2593), .Y(dp.rf._abc_6362_n3194) );
	NAND2X1 NAND2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2595) );
	NAND2X1 NAND2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<5>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2596) );
	NAND2X1 NAND2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2595), .B(dp.rf._abc_6362_n2596), .Y(dp.rf._abc_6362_n3195) );
	NAND2X1 NAND2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2598) );
	NAND2X1 NAND2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<6>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2599) );
	NAND2X1 NAND2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2598), .B(dp.rf._abc_6362_n2599), .Y(dp.rf._abc_6362_n3196) );
	NAND2X1 NAND2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2601) );
	NAND2X1 NAND2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<7>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2602) );
	NAND2X1 NAND2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2601), .B(dp.rf._abc_6362_n2602), .Y(dp.rf._abc_6362_n3197) );
	NAND2X1 NAND2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2604) );
	NAND2X1 NAND2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<8>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2605) );
	NAND2X1 NAND2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2604), .B(dp.rf._abc_6362_n2605), .Y(dp.rf._abc_6362_n3198) );
	NAND2X1 NAND2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2607) );
	NAND2X1 NAND2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<9>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2608) );
	NAND2X1 NAND2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2607), .B(dp.rf._abc_6362_n2608), .Y(dp.rf._abc_6362_n3199) );
	NAND2X1 NAND2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2610) );
	NAND2X1 NAND2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<10>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2611) );
	NAND2X1 NAND2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2610), .B(dp.rf._abc_6362_n2611), .Y(dp.rf._abc_6362_n3200) );
	NAND2X1 NAND2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2613) );
	NAND2X1 NAND2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<11>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2614) );
	NAND2X1 NAND2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2613), .B(dp.rf._abc_6362_n2614), .Y(dp.rf._abc_6362_n3201) );
	NAND2X1 NAND2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2616) );
	NAND2X1 NAND2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<12>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2617) );
	NAND2X1 NAND2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2616), .B(dp.rf._abc_6362_n2617), .Y(dp.rf._abc_6362_n3202) );
	NAND2X1 NAND2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2619) );
	NAND2X1 NAND2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<13>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2620) );
	NAND2X1 NAND2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2619), .B(dp.rf._abc_6362_n2620), .Y(dp.rf._abc_6362_n3203) );
	NAND2X1 NAND2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2622) );
	NAND2X1 NAND2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<14>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2623) );
	NAND2X1 NAND2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2622), .B(dp.rf._abc_6362_n2623), .Y(dp.rf._abc_6362_n3204) );
	NAND2X1 NAND2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2625) );
	NAND2X1 NAND2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<15>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2626) );
	NAND2X1 NAND2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2625), .B(dp.rf._abc_6362_n2626), .Y(dp.rf._abc_6362_n3205) );
	NAND2X1 NAND2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2628) );
	NAND2X1 NAND2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<16>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2629) );
	NAND2X1 NAND2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2628), .B(dp.rf._abc_6362_n2629), .Y(dp.rf._abc_6362_n3206) );
	NAND2X1 NAND2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2631) );
	NAND2X1 NAND2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<17>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2632) );
	NAND2X1 NAND2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2631), .B(dp.rf._abc_6362_n2632), .Y(dp.rf._abc_6362_n3207) );
	NAND2X1 NAND2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2634) );
	NAND2X1 NAND2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<18>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2635) );
	NAND2X1 NAND2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2634), .B(dp.rf._abc_6362_n2635), .Y(dp.rf._abc_6362_n3208) );
	NAND2X1 NAND2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2637) );
	NAND2X1 NAND2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<19>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2638) );
	NAND2X1 NAND2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2637), .B(dp.rf._abc_6362_n2638), .Y(dp.rf._abc_6362_n3209) );
	NAND2X1 NAND2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2640) );
	NAND2X1 NAND2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<20>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2641) );
	NAND2X1 NAND2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2640), .B(dp.rf._abc_6362_n2641), .Y(dp.rf._abc_6362_n3210) );
	NAND2X1 NAND2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2643) );
	NAND2X1 NAND2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<21>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2644) );
	NAND2X1 NAND2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2643), .B(dp.rf._abc_6362_n2644), .Y(dp.rf._abc_6362_n3211) );
	NAND2X1 NAND2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2646) );
	NAND2X1 NAND2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<22>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2647) );
	NAND2X1 NAND2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2646), .B(dp.rf._abc_6362_n2647), .Y(dp.rf._abc_6362_n3212) );
	NAND2X1 NAND2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2649) );
	NAND2X1 NAND2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<23>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2650) );
	NAND2X1 NAND2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2649), .B(dp.rf._abc_6362_n2650), .Y(dp.rf._abc_6362_n3213) );
	NAND2X1 NAND2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2652) );
	NAND2X1 NAND2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<24>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2653) );
	NAND2X1 NAND2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2652), .B(dp.rf._abc_6362_n2653), .Y(dp.rf._abc_6362_n3214) );
	NAND2X1 NAND2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2655) );
	NAND2X1 NAND2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<25>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2656) );
	NAND2X1 NAND2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2655), .B(dp.rf._abc_6362_n2656), .Y(dp.rf._abc_6362_n3215) );
	NAND2X1 NAND2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2658) );
	NAND2X1 NAND2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<26>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2659) );
	NAND2X1 NAND2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2658), .B(dp.rf._abc_6362_n2659), .Y(dp.rf._abc_6362_n3216) );
	NAND2X1 NAND2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2661) );
	NAND2X1 NAND2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<27>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2662) );
	NAND2X1 NAND2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2661), .B(dp.rf._abc_6362_n2662), .Y(dp.rf._abc_6362_n3217) );
	NAND2X1 NAND2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2664) );
	NAND2X1 NAND2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<28>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2665) );
	NAND2X1 NAND2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2664), .B(dp.rf._abc_6362_n2665), .Y(dp.rf._abc_6362_n3218) );
	NAND2X1 NAND2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2667) );
	NAND2X1 NAND2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<29>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2668) );
	NAND2X1 NAND2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2667), .B(dp.rf._abc_6362_n2668), .Y(dp.rf._abc_6362_n3219) );
	NAND2X1 NAND2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2670) );
	NAND2X1 NAND2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<30>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2671) );
	NAND2X1 NAND2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2670), .B(dp.rf._abc_6362_n2671), .Y(dp.rf._abc_6362_n3220) );
	NAND2X1 NAND2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n2578), .Y(dp.rf._abc_6362_n2673) );
	NAND2X1 NAND2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_13_<31>), .B(dp.rf._abc_6362_n2580), .Y(dp.rf._abc_6362_n2674) );
	NAND2X1 NAND2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2673), .B(dp.rf._abc_6362_n2674), .Y(dp.rf._abc_6362_n3221) );
	NAND2X1 NAND2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2273), .B(dp.rf._abc_6362_n2476), .Y(dp.rf._abc_6362_n2676) );
	NOR2X1 NOR2X1_196 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n2676), .Y(dp.rf._abc_6362_n2677) );
	NAND2X1 NAND2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2678) );
	INVX8 INVX8_10 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2679) );
	NAND2X1 NAND2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<0>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2680) );
	NAND2X1 NAND2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2678), .B(dp.rf._abc_6362_n2680), .Y(dp.rf._abc_6362_n3222) );
	NAND2X1 NAND2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2682) );
	NAND2X1 NAND2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<1>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2683) );
	NAND2X1 NAND2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2682), .B(dp.rf._abc_6362_n2683), .Y(dp.rf._abc_6362_n3223) );
	NAND2X1 NAND2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2685) );
	NAND2X1 NAND2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<2>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2686) );
	NAND2X1 NAND2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2685), .B(dp.rf._abc_6362_n2686), .Y(dp.rf._abc_6362_n3224) );
	NAND2X1 NAND2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2688) );
	NAND2X1 NAND2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<3>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2689) );
	NAND2X1 NAND2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2688), .B(dp.rf._abc_6362_n2689), .Y(dp.rf._abc_6362_n3225) );
	NAND2X1 NAND2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2691) );
	NAND2X1 NAND2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<4>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2692) );
	NAND2X1 NAND2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2691), .B(dp.rf._abc_6362_n2692), .Y(dp.rf._abc_6362_n3226) );
	NAND2X1 NAND2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2694) );
	NAND2X1 NAND2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<5>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2695) );
	NAND2X1 NAND2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2694), .B(dp.rf._abc_6362_n2695), .Y(dp.rf._abc_6362_n3227) );
	NAND2X1 NAND2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2697) );
	NAND2X1 NAND2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<6>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2698) );
	NAND2X1 NAND2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2697), .B(dp.rf._abc_6362_n2698), .Y(dp.rf._abc_6362_n3228) );
	NAND2X1 NAND2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2700) );
	NAND2X1 NAND2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<7>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2701) );
	NAND2X1 NAND2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2700), .B(dp.rf._abc_6362_n2701), .Y(dp.rf._abc_6362_n3229) );
	NAND2X1 NAND2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2703) );
	NAND2X1 NAND2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<8>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2704) );
	NAND2X1 NAND2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2703), .B(dp.rf._abc_6362_n2704), .Y(dp.rf._abc_6362_n3230) );
	NAND2X1 NAND2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2706) );
	NAND2X1 NAND2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<9>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2707) );
	NAND2X1 NAND2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2706), .B(dp.rf._abc_6362_n2707), .Y(dp.rf._abc_6362_n3231) );
	NAND2X1 NAND2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2709) );
	NAND2X1 NAND2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<10>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2710) );
	NAND2X1 NAND2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2709), .B(dp.rf._abc_6362_n2710), .Y(dp.rf._abc_6362_n3232) );
	NAND2X1 NAND2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2712) );
	NAND2X1 NAND2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<11>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2713) );
	NAND2X1 NAND2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2712), .B(dp.rf._abc_6362_n2713), .Y(dp.rf._abc_6362_n3233) );
	NAND2X1 NAND2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2715) );
	NAND2X1 NAND2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<12>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2716) );
	NAND2X1 NAND2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2715), .B(dp.rf._abc_6362_n2716), .Y(dp.rf._abc_6362_n3234) );
	NAND2X1 NAND2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2718) );
	NAND2X1 NAND2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<13>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2719) );
	NAND2X1 NAND2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2718), .B(dp.rf._abc_6362_n2719), .Y(dp.rf._abc_6362_n3235) );
	NAND2X1 NAND2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2721) );
	NAND2X1 NAND2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<14>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2722) );
	NAND2X1 NAND2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2721), .B(dp.rf._abc_6362_n2722), .Y(dp.rf._abc_6362_n3236) );
	NAND2X1 NAND2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2724) );
	NAND2X1 NAND2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<15>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2725) );
	NAND2X1 NAND2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2724), .B(dp.rf._abc_6362_n2725), .Y(dp.rf._abc_6362_n3237) );
	NAND2X1 NAND2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2727) );
	NAND2X1 NAND2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<16>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2728) );
	NAND2X1 NAND2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2727), .B(dp.rf._abc_6362_n2728), .Y(dp.rf._abc_6362_n3238) );
	NAND2X1 NAND2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2730) );
	NAND2X1 NAND2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<17>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2731) );
	NAND2X1 NAND2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2730), .B(dp.rf._abc_6362_n2731), .Y(dp.rf._abc_6362_n3239) );
	NAND2X1 NAND2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2733) );
	NAND2X1 NAND2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<18>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2734) );
	NAND2X1 NAND2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2733), .B(dp.rf._abc_6362_n2734), .Y(dp.rf._abc_6362_n3240) );
	NAND2X1 NAND2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2736) );
	NAND2X1 NAND2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<19>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2737) );
	NAND2X1 NAND2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2736), .B(dp.rf._abc_6362_n2737), .Y(dp.rf._abc_6362_n3241) );
	NAND2X1 NAND2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2739) );
	NAND2X1 NAND2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<20>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2740) );
	NAND2X1 NAND2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2739), .B(dp.rf._abc_6362_n2740), .Y(dp.rf._abc_6362_n3242) );
	NAND2X1 NAND2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2742) );
	NAND2X1 NAND2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<21>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2743) );
	NAND2X1 NAND2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2742), .B(dp.rf._abc_6362_n2743), .Y(dp.rf._abc_6362_n3243) );
	NAND2X1 NAND2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2745) );
	NAND2X1 NAND2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<22>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2746) );
	NAND2X1 NAND2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2745), .B(dp.rf._abc_6362_n2746), .Y(dp.rf._abc_6362_n3244) );
	NAND2X1 NAND2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2748) );
	NAND2X1 NAND2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<23>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2749) );
	NAND2X1 NAND2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2748), .B(dp.rf._abc_6362_n2749), .Y(dp.rf._abc_6362_n3245) );
	NAND2X1 NAND2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2751) );
	NAND2X1 NAND2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<24>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2752) );
	NAND2X1 NAND2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2751), .B(dp.rf._abc_6362_n2752), .Y(dp.rf._abc_6362_n3246) );
	NAND2X1 NAND2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2754) );
	NAND2X1 NAND2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<25>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2755) );
	NAND2X1 NAND2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2754), .B(dp.rf._abc_6362_n2755), .Y(dp.rf._abc_6362_n3247) );
	NAND2X1 NAND2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2757) );
	NAND2X1 NAND2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<26>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2758) );
	NAND2X1 NAND2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2757), .B(dp.rf._abc_6362_n2758), .Y(dp.rf._abc_6362_n3248) );
	NAND2X1 NAND2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2760) );
	NAND2X1 NAND2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<27>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2761) );
	NAND2X1 NAND2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2760), .B(dp.rf._abc_6362_n2761), .Y(dp.rf._abc_6362_n3249) );
	NAND2X1 NAND2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2763) );
	NAND2X1 NAND2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<28>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2764) );
	NAND2X1 NAND2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2763), .B(dp.rf._abc_6362_n2764), .Y(dp.rf._abc_6362_n3250) );
	NAND2X1 NAND2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2766) );
	NAND2X1 NAND2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<29>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2767) );
	NAND2X1 NAND2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2766), .B(dp.rf._abc_6362_n2767), .Y(dp.rf._abc_6362_n3251) );
	NAND2X1 NAND2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2769) );
	NAND2X1 NAND2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<30>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2770) );
	NAND2X1 NAND2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2769), .B(dp.rf._abc_6362_n2770), .Y(dp.rf._abc_6362_n3252) );
	NAND2X1 NAND2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n2677), .Y(dp.rf._abc_6362_n2772) );
	NAND2X1 NAND2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<31>), .B(dp.rf._abc_6362_n2679), .Y(dp.rf._abc_6362_n2773) );
	NAND2X1 NAND2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2772), .B(dp.rf._abc_6362_n2773), .Y(dp.rf._abc_6362_n3253) );
	NAND2X1 NAND2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2376), .B(dp.rf._abc_6362_n2476), .Y(dp.rf._abc_6362_n2775) );
	NOR2X1 NOR2X1_197 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n2775), .Y(dp.rf._abc_6362_n2776) );
	NAND2X1 NAND2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2777) );
	INVX8 INVX8_11 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2778) );
	NAND2X1 NAND2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<0>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2779) );
	NAND2X1 NAND2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2777), .B(dp.rf._abc_6362_n2779), .Y(dp.rf._abc_6362_n3254) );
	NAND2X1 NAND2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2781) );
	NAND2X1 NAND2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<1>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2782) );
	NAND2X1 NAND2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2781), .B(dp.rf._abc_6362_n2782), .Y(dp.rf._abc_6362_n3255) );
	NAND2X1 NAND2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2784) );
	NAND2X1 NAND2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<2>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2785) );
	NAND2X1 NAND2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2784), .B(dp.rf._abc_6362_n2785), .Y(dp.rf._abc_6362_n3256) );
	NAND2X1 NAND2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2787) );
	NAND2X1 NAND2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<3>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2788) );
	NAND2X1 NAND2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2787), .B(dp.rf._abc_6362_n2788), .Y(dp.rf._abc_6362_n3257) );
	NAND2X1 NAND2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2790) );
	NAND2X1 NAND2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<4>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2791) );
	NAND2X1 NAND2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2790), .B(dp.rf._abc_6362_n2791), .Y(dp.rf._abc_6362_n3258) );
	NAND2X1 NAND2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2793) );
	NAND2X1 NAND2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<5>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2794) );
	NAND2X1 NAND2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2793), .B(dp.rf._abc_6362_n2794), .Y(dp.rf._abc_6362_n3259) );
	NAND2X1 NAND2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2796) );
	NAND2X1 NAND2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<6>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2797) );
	NAND2X1 NAND2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2796), .B(dp.rf._abc_6362_n2797), .Y(dp.rf._abc_6362_n3260) );
	NAND2X1 NAND2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2799) );
	NAND2X1 NAND2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<7>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2800) );
	NAND2X1 NAND2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2799), .B(dp.rf._abc_6362_n2800), .Y(dp.rf._abc_6362_n3261) );
	NAND2X1 NAND2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2802) );
	NAND2X1 NAND2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<8>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2803) );
	NAND2X1 NAND2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2802), .B(dp.rf._abc_6362_n2803), .Y(dp.rf._abc_6362_n3262) );
	NAND2X1 NAND2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2805) );
	NAND2X1 NAND2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<9>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2806) );
	NAND2X1 NAND2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2805), .B(dp.rf._abc_6362_n2806), .Y(dp.rf._abc_6362_n3263) );
	NAND2X1 NAND2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2808) );
	NAND2X1 NAND2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<10>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2809) );
	NAND2X1 NAND2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2808), .B(dp.rf._abc_6362_n2809), .Y(dp.rf._abc_6362_n3264) );
	NAND2X1 NAND2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2811) );
	NAND2X1 NAND2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<11>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2812) );
	NAND2X1 NAND2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2811), .B(dp.rf._abc_6362_n2812), .Y(dp.rf._abc_6362_n3265) );
	NAND2X1 NAND2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2814) );
	NAND2X1 NAND2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<12>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2815) );
	NAND2X1 NAND2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2814), .B(dp.rf._abc_6362_n2815), .Y(dp.rf._abc_6362_n3266) );
	NAND2X1 NAND2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2817) );
	NAND2X1 NAND2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<13>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2818) );
	NAND2X1 NAND2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2817), .B(dp.rf._abc_6362_n2818), .Y(dp.rf._abc_6362_n3267) );
	NAND2X1 NAND2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2820) );
	NAND2X1 NAND2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<14>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2821) );
	NAND2X1 NAND2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2820), .B(dp.rf._abc_6362_n2821), .Y(dp.rf._abc_6362_n3268) );
	NAND2X1 NAND2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2823) );
	NAND2X1 NAND2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<15>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2824) );
	NAND2X1 NAND2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2823), .B(dp.rf._abc_6362_n2824), .Y(dp.rf._abc_6362_n3269) );
	NAND2X1 NAND2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2826) );
	NAND2X1 NAND2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<16>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2827) );
	NAND2X1 NAND2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2826), .B(dp.rf._abc_6362_n2827), .Y(dp.rf._abc_6362_n3270) );
	NAND2X1 NAND2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2829) );
	NAND2X1 NAND2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<17>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2830) );
	NAND2X1 NAND2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2829), .B(dp.rf._abc_6362_n2830), .Y(dp.rf._abc_6362_n3271) );
	NAND2X1 NAND2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2832) );
	NAND2X1 NAND2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<18>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2833) );
	NAND2X1 NAND2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2832), .B(dp.rf._abc_6362_n2833), .Y(dp.rf._abc_6362_n3272) );
	NAND2X1 NAND2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2835) );
	NAND2X1 NAND2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<19>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2836) );
	NAND2X1 NAND2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2835), .B(dp.rf._abc_6362_n2836), .Y(dp.rf._abc_6362_n3273) );
	NAND2X1 NAND2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2838) );
	NAND2X1 NAND2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<20>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2839) );
	NAND2X1 NAND2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2838), .B(dp.rf._abc_6362_n2839), .Y(dp.rf._abc_6362_n3274) );
	NAND2X1 NAND2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2841) );
	NAND2X1 NAND2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<21>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2842) );
	NAND2X1 NAND2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2841), .B(dp.rf._abc_6362_n2842), .Y(dp.rf._abc_6362_n3275) );
	NAND2X1 NAND2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2844) );
	NAND2X1 NAND2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<22>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2845) );
	NAND2X1 NAND2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2844), .B(dp.rf._abc_6362_n2845), .Y(dp.rf._abc_6362_n3276) );
	NAND2X1 NAND2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2847) );
	NAND2X1 NAND2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<23>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2848) );
	NAND2X1 NAND2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2847), .B(dp.rf._abc_6362_n2848), .Y(dp.rf._abc_6362_n3277) );
	NAND2X1 NAND2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2850) );
	NAND2X1 NAND2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<24>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2851) );
	NAND2X1 NAND2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2850), .B(dp.rf._abc_6362_n2851), .Y(dp.rf._abc_6362_n3278) );
	NAND2X1 NAND2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2853) );
	NAND2X1 NAND2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<25>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2854) );
	NAND2X1 NAND2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2853), .B(dp.rf._abc_6362_n2854), .Y(dp.rf._abc_6362_n3279) );
	NAND2X1 NAND2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2856) );
	NAND2X1 NAND2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<26>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2857) );
	NAND2X1 NAND2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2856), .B(dp.rf._abc_6362_n2857), .Y(dp.rf._abc_6362_n3280) );
	NAND2X1 NAND2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2859) );
	NAND2X1 NAND2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<27>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2860) );
	NAND2X1 NAND2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2859), .B(dp.rf._abc_6362_n2860), .Y(dp.rf._abc_6362_n3281) );
	NAND2X1 NAND2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2862) );
	NAND2X1 NAND2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<28>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2863) );
	NAND2X1 NAND2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2862), .B(dp.rf._abc_6362_n2863), .Y(dp.rf._abc_6362_n3282) );
	NAND2X1 NAND2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2865) );
	NAND2X1 NAND2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<29>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2866) );
	NAND2X1 NAND2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2865), .B(dp.rf._abc_6362_n2866), .Y(dp.rf._abc_6362_n3283) );
	NAND2X1 NAND2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2868) );
	NAND2X1 NAND2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<30>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2869) );
	NAND2X1 NAND2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2868), .B(dp.rf._abc_6362_n2869), .Y(dp.rf._abc_6362_n3284) );
	NAND2X1 NAND2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n2776), .Y(dp.rf._abc_6362_n2871) );
	NAND2X1 NAND2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_15_<31>), .B(dp.rf._abc_6362_n2778), .Y(dp.rf._abc_6362_n2872) );
	NAND2X1 NAND2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2871), .B(dp.rf._abc_6362_n2872), .Y(dp.rf._abc_6362_n3285) );
	AND2X2 AND2X2_75 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_8_), .B(dp.writereg_4_), .Y(dp.rf._abc_6362_n2874) );
	INVX4 INVX4_3 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2874), .Y(dp.rf._abc_6362_n2875) );
	NOR2X1 NOR2X1_198 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n2173), .Y(dp.rf._abc_6362_n2876) );
	NAND2X1 NAND2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2877) );
	INVX8 INVX8_12 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2878) );
	NAND2X1 NAND2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<0>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2879) );
	NAND2X1 NAND2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2877), .B(dp.rf._abc_6362_n2879), .Y(dp.rf._abc_6362_n3286) );
	NAND2X1 NAND2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2881) );
	NAND2X1 NAND2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<1>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2882) );
	NAND2X1 NAND2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2881), .B(dp.rf._abc_6362_n2882), .Y(dp.rf._abc_6362_n3287) );
	NAND2X1 NAND2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2884) );
	NAND2X1 NAND2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<2>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2885) );
	NAND2X1 NAND2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2884), .B(dp.rf._abc_6362_n2885), .Y(dp.rf._abc_6362_n3288) );
	NAND2X1 NAND2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2887) );
	NAND2X1 NAND2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<3>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2888) );
	NAND2X1 NAND2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2887), .B(dp.rf._abc_6362_n2888), .Y(dp.rf._abc_6362_n3289) );
	NAND2X1 NAND2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2890) );
	NAND2X1 NAND2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<4>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2891) );
	NAND2X1 NAND2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2890), .B(dp.rf._abc_6362_n2891), .Y(dp.rf._abc_6362_n3290) );
	NAND2X1 NAND2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2893) );
	NAND2X1 NAND2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<5>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2894) );
	NAND2X1 NAND2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2893), .B(dp.rf._abc_6362_n2894), .Y(dp.rf._abc_6362_n3291) );
	NAND2X1 NAND2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2896) );
	NAND2X1 NAND2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<6>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2897) );
	NAND2X1 NAND2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2896), .B(dp.rf._abc_6362_n2897), .Y(dp.rf._abc_6362_n3292) );
	NAND2X1 NAND2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2899) );
	NAND2X1 NAND2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<7>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2900) );
	NAND2X1 NAND2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2899), .B(dp.rf._abc_6362_n2900), .Y(dp.rf._abc_6362_n3293) );
	NAND2X1 NAND2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2902) );
	NAND2X1 NAND2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<8>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2903) );
	NAND2X1 NAND2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2902), .B(dp.rf._abc_6362_n2903), .Y(dp.rf._abc_6362_n3294) );
	NAND2X1 NAND2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2905) );
	NAND2X1 NAND2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<9>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2906) );
	NAND2X1 NAND2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2905), .B(dp.rf._abc_6362_n2906), .Y(dp.rf._abc_6362_n3295) );
	NAND2X1 NAND2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2908) );
	NAND2X1 NAND2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<10>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2909) );
	NAND2X1 NAND2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2908), .B(dp.rf._abc_6362_n2909), .Y(dp.rf._abc_6362_n3296) );
	NAND2X1 NAND2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2911) );
	NAND2X1 NAND2X1_1403 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<11>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2912) );
	NAND2X1 NAND2X1_1404 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2911), .B(dp.rf._abc_6362_n2912), .Y(dp.rf._abc_6362_n3297) );
	NAND2X1 NAND2X1_1405 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2914) );
	NAND2X1 NAND2X1_1406 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<12>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2915) );
	NAND2X1 NAND2X1_1407 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2914), .B(dp.rf._abc_6362_n2915), .Y(dp.rf._abc_6362_n3298) );
	NAND2X1 NAND2X1_1408 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2917) );
	NAND2X1 NAND2X1_1409 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<13>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2918) );
	NAND2X1 NAND2X1_1410 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2917), .B(dp.rf._abc_6362_n2918), .Y(dp.rf._abc_6362_n3299) );
	NAND2X1 NAND2X1_1411 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2920) );
	NAND2X1 NAND2X1_1412 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<14>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2921) );
	NAND2X1 NAND2X1_1413 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2920), .B(dp.rf._abc_6362_n2921), .Y(dp.rf._abc_6362_n3300) );
	NAND2X1 NAND2X1_1414 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2923) );
	NAND2X1 NAND2X1_1415 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<15>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2924) );
	NAND2X1 NAND2X1_1416 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2923), .B(dp.rf._abc_6362_n2924), .Y(dp.rf._abc_6362_n3301) );
	NAND2X1 NAND2X1_1417 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2926) );
	NAND2X1 NAND2X1_1418 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<16>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2927) );
	NAND2X1 NAND2X1_1419 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2926), .B(dp.rf._abc_6362_n2927), .Y(dp.rf._abc_6362_n3302) );
	NAND2X1 NAND2X1_1420 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2929) );
	NAND2X1 NAND2X1_1421 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<17>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2930) );
	NAND2X1 NAND2X1_1422 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2929), .B(dp.rf._abc_6362_n2930), .Y(dp.rf._abc_6362_n3303) );
	NAND2X1 NAND2X1_1423 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2932) );
	NAND2X1 NAND2X1_1424 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<18>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2933) );
	NAND2X1 NAND2X1_1425 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2932), .B(dp.rf._abc_6362_n2933), .Y(dp.rf._abc_6362_n3304) );
	NAND2X1 NAND2X1_1426 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2935) );
	NAND2X1 NAND2X1_1427 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<19>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2936) );
	NAND2X1 NAND2X1_1428 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2935), .B(dp.rf._abc_6362_n2936), .Y(dp.rf._abc_6362_n3305) );
	NAND2X1 NAND2X1_1429 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2938) );
	NAND2X1 NAND2X1_1430 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<20>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2939) );
	NAND2X1 NAND2X1_1431 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2938), .B(dp.rf._abc_6362_n2939), .Y(dp.rf._abc_6362_n3306) );
	NAND2X1 NAND2X1_1432 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2941) );
	NAND2X1 NAND2X1_1433 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<21>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2942) );
	NAND2X1 NAND2X1_1434 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2941), .B(dp.rf._abc_6362_n2942), .Y(dp.rf._abc_6362_n3307) );
	NAND2X1 NAND2X1_1435 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2944) );
	NAND2X1 NAND2X1_1436 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<22>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2945) );
	NAND2X1 NAND2X1_1437 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2944), .B(dp.rf._abc_6362_n2945), .Y(dp.rf._abc_6362_n3308) );
	NAND2X1 NAND2X1_1438 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2947) );
	NAND2X1 NAND2X1_1439 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<23>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2948) );
	NAND2X1 NAND2X1_1440 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2947), .B(dp.rf._abc_6362_n2948), .Y(dp.rf._abc_6362_n3309) );
	NAND2X1 NAND2X1_1441 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2950) );
	NAND2X1 NAND2X1_1442 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<24>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2951) );
	NAND2X1 NAND2X1_1443 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2950), .B(dp.rf._abc_6362_n2951), .Y(dp.rf._abc_6362_n3310) );
	NAND2X1 NAND2X1_1444 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2953) );
	NAND2X1 NAND2X1_1445 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<25>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2954) );
	NAND2X1 NAND2X1_1446 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2953), .B(dp.rf._abc_6362_n2954), .Y(dp.rf._abc_6362_n3311) );
	NAND2X1 NAND2X1_1447 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2956) );
	NAND2X1 NAND2X1_1448 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<26>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2957) );
	NAND2X1 NAND2X1_1449 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2956), .B(dp.rf._abc_6362_n2957), .Y(dp.rf._abc_6362_n3312) );
	NAND2X1 NAND2X1_1450 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2959) );
	NAND2X1 NAND2X1_1451 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<27>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2960) );
	NAND2X1 NAND2X1_1452 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2959), .B(dp.rf._abc_6362_n2960), .Y(dp.rf._abc_6362_n3313) );
	NAND2X1 NAND2X1_1453 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2962) );
	NAND2X1 NAND2X1_1454 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<28>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2963) );
	NAND2X1 NAND2X1_1455 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2962), .B(dp.rf._abc_6362_n2963), .Y(dp.rf._abc_6362_n3314) );
	NAND2X1 NAND2X1_1456 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2965) );
	NAND2X1 NAND2X1_1457 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<29>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2966) );
	NAND2X1 NAND2X1_1458 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2965), .B(dp.rf._abc_6362_n2966), .Y(dp.rf._abc_6362_n3315) );
	NAND2X1 NAND2X1_1459 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2968) );
	NAND2X1 NAND2X1_1460 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<30>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2969) );
	NAND2X1 NAND2X1_1461 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2968), .B(dp.rf._abc_6362_n2969), .Y(dp.rf._abc_6362_n3316) );
	NAND2X1 NAND2X1_1462 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n2876), .Y(dp.rf._abc_6362_n2971) );
	NAND2X1 NAND2X1_1463 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<31>), .B(dp.rf._abc_6362_n2878), .Y(dp.rf._abc_6362_n2972) );
	NAND2X1 NAND2X1_1464 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2971), .B(dp.rf._abc_6362_n2972), .Y(dp.rf._abc_6362_n3317) );
	NAND2X1 NAND2X1_1465 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2172), .B(dp.rf._abc_6362_n2576), .Y(dp.rf._abc_6362_n2974) );
	NOR2X1 NOR2X1_199 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n2974), .Y(dp.rf._abc_6362_n2975) );
	NAND2X1 NAND2X1_1466 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n2976) );
	INVX8 INVX8_13 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n2977) );
	NAND2X1 NAND2X1_1467 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<0>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n2978) );
	NAND2X1 NAND2X1_1468 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2976), .B(dp.rf._abc_6362_n2978), .Y(dp.rf._abc_6362_n3318) );
	NAND2X1 NAND2X1_1469 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n2980) );
	NAND2X1 NAND2X1_1470 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<1>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n2981) );
	NAND2X1 NAND2X1_1471 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2980), .B(dp.rf._abc_6362_n2981), .Y(dp.rf._abc_6362_n3319) );
	NAND2X1 NAND2X1_1472 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n2983) );
	NAND2X1 NAND2X1_1473 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<2>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n2984) );
	NAND2X1 NAND2X1_1474 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2983), .B(dp.rf._abc_6362_n2984), .Y(dp.rf._abc_6362_n3320) );
	NAND2X1 NAND2X1_1475 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n2986) );
	NAND2X1 NAND2X1_1476 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<3>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n2987) );
	NAND2X1 NAND2X1_1477 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2986), .B(dp.rf._abc_6362_n2987), .Y(dp.rf._abc_6362_n3321) );
	NAND2X1 NAND2X1_1478 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n2989) );
	NAND2X1 NAND2X1_1479 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<4>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n2990) );
	NAND2X1 NAND2X1_1480 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2989), .B(dp.rf._abc_6362_n2990), .Y(dp.rf._abc_6362_n3322) );
	NAND2X1 NAND2X1_1481 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n2992) );
	NAND2X1 NAND2X1_1482 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<5>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n2993) );
	NAND2X1 NAND2X1_1483 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2992), .B(dp.rf._abc_6362_n2993), .Y(dp.rf._abc_6362_n3323) );
	NAND2X1 NAND2X1_1484 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n2995) );
	NAND2X1 NAND2X1_1485 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<6>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n2996) );
	NAND2X1 NAND2X1_1486 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2995), .B(dp.rf._abc_6362_n2996), .Y(dp.rf._abc_6362_n3324) );
	NAND2X1 NAND2X1_1487 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n2998) );
	NAND2X1 NAND2X1_1488 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<7>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n2999) );
	NAND2X1 NAND2X1_1489 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2998), .B(dp.rf._abc_6362_n2999), .Y(dp.rf._abc_6362_n3325) );
	NAND2X1 NAND2X1_1490 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3001) );
	NAND2X1 NAND2X1_1491 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<8>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3002) );
	NAND2X1 NAND2X1_1492 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3001), .B(dp.rf._abc_6362_n3002), .Y(dp.rf._abc_6362_n3326) );
	NAND2X1 NAND2X1_1493 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3004) );
	NAND2X1 NAND2X1_1494 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<9>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3005) );
	NAND2X1 NAND2X1_1495 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3004), .B(dp.rf._abc_6362_n3005), .Y(dp.rf._abc_6362_n3327) );
	NAND2X1 NAND2X1_1496 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3007) );
	NAND2X1 NAND2X1_1497 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<10>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3008) );
	NAND2X1 NAND2X1_1498 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3007), .B(dp.rf._abc_6362_n3008), .Y(dp.rf._abc_6362_n3328) );
	NAND2X1 NAND2X1_1499 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3010) );
	NAND2X1 NAND2X1_1500 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<11>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3011) );
	NAND2X1 NAND2X1_1501 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3010), .B(dp.rf._abc_6362_n3011), .Y(dp.rf._abc_6362_n3329) );
	NAND2X1 NAND2X1_1502 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3013) );
	NAND2X1 NAND2X1_1503 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<12>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3014) );
	NAND2X1 NAND2X1_1504 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3013), .B(dp.rf._abc_6362_n3014), .Y(dp.rf._abc_6362_n3330) );
	NAND2X1 NAND2X1_1505 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3016) );
	NAND2X1 NAND2X1_1506 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<13>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3017) );
	NAND2X1 NAND2X1_1507 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3016), .B(dp.rf._abc_6362_n3017), .Y(dp.rf._abc_6362_n3331) );
	NAND2X1 NAND2X1_1508 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3019) );
	NAND2X1 NAND2X1_1509 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<14>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3020) );
	NAND2X1 NAND2X1_1510 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3019), .B(dp.rf._abc_6362_n3020), .Y(dp.rf._abc_6362_n3332) );
	NAND2X1 NAND2X1_1511 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3022) );
	NAND2X1 NAND2X1_1512 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<15>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3023) );
	NAND2X1 NAND2X1_1513 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3022), .B(dp.rf._abc_6362_n3023), .Y(dp.rf._abc_6362_n3333) );
	NAND2X1 NAND2X1_1514 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3025) );
	NAND2X1 NAND2X1_1515 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<16>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3026) );
	NAND2X1 NAND2X1_1516 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3025), .B(dp.rf._abc_6362_n3026), .Y(dp.rf._abc_6362_n3334) );
	NAND2X1 NAND2X1_1517 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3028) );
	NAND2X1 NAND2X1_1518 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<17>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3029) );
	NAND2X1 NAND2X1_1519 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3028), .B(dp.rf._abc_6362_n3029), .Y(dp.rf._abc_6362_n3335) );
	NAND2X1 NAND2X1_1520 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3031_1) );
	NAND2X1 NAND2X1_1521 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<18>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3032) );
	NAND2X1 NAND2X1_1522 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3031_1), .B(dp.rf._abc_6362_n3032), .Y(dp.rf._abc_6362_n3336) );
	NAND2X1 NAND2X1_1523 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3034) );
	NAND2X1 NAND2X1_1524 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<19>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3035_1) );
	NAND2X1 NAND2X1_1525 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3034), .B(dp.rf._abc_6362_n3035_1), .Y(dp.rf._abc_6362_n3337) );
	NAND2X1 NAND2X1_1526 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3037_1) );
	NAND2X1 NAND2X1_1527 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<20>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3038) );
	NAND2X1 NAND2X1_1528 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3037_1), .B(dp.rf._abc_6362_n3038), .Y(dp.rf._abc_6362_n3338) );
	NAND2X1 NAND2X1_1529 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3040) );
	NAND2X1 NAND2X1_1530 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<21>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3041_1) );
	NAND2X1 NAND2X1_1531 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3040), .B(dp.rf._abc_6362_n3041_1), .Y(dp.rf._abc_6362_n3339) );
	NAND2X1 NAND2X1_1532 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3043_1) );
	NAND2X1 NAND2X1_1533 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<22>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3044) );
	NAND2X1 NAND2X1_1534 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3043_1), .B(dp.rf._abc_6362_n3044), .Y(dp.rf._abc_6362_n3340) );
	NAND2X1 NAND2X1_1535 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3046) );
	NAND2X1 NAND2X1_1536 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<23>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3047_1) );
	NAND2X1 NAND2X1_1537 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3046), .B(dp.rf._abc_6362_n3047_1), .Y(dp.rf._abc_6362_n3341) );
	NAND2X1 NAND2X1_1538 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3049_1) );
	NAND2X1 NAND2X1_1539 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<24>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3050) );
	NAND2X1 NAND2X1_1540 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3049_1), .B(dp.rf._abc_6362_n3050), .Y(dp.rf._abc_6362_n3342) );
	NAND2X1 NAND2X1_1541 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3052) );
	NAND2X1 NAND2X1_1542 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<25>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3053_1) );
	NAND2X1 NAND2X1_1543 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3052), .B(dp.rf._abc_6362_n3053_1), .Y(dp.rf._abc_6362_n3343) );
	NAND2X1 NAND2X1_1544 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3055_1) );
	NAND2X1 NAND2X1_1545 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<26>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3056) );
	NAND2X1 NAND2X1_1546 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3055_1), .B(dp.rf._abc_6362_n3056), .Y(dp.rf._abc_6362_n3344) );
	NAND2X1 NAND2X1_1547 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3058) );
	NAND2X1 NAND2X1_1548 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<27>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3059_1) );
	NAND2X1 NAND2X1_1549 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3058), .B(dp.rf._abc_6362_n3059_1), .Y(dp.rf._abc_6362_n3345) );
	NAND2X1 NAND2X1_1550 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3061_1) );
	NAND2X1 NAND2X1_1551 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<28>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3062) );
	NAND2X1 NAND2X1_1552 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3061_1), .B(dp.rf._abc_6362_n3062), .Y(dp.rf._abc_6362_n3346) );
	NAND2X1 NAND2X1_1553 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3064) );
	NAND2X1 NAND2X1_1554 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<29>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3065_1) );
	NAND2X1 NAND2X1_1555 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3064), .B(dp.rf._abc_6362_n3065_1), .Y(dp.rf._abc_6362_n3347) );
	NAND2X1 NAND2X1_1556 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3067_1) );
	NAND2X1 NAND2X1_1557 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<30>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3068) );
	NAND2X1 NAND2X1_1558 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3067_1), .B(dp.rf._abc_6362_n3068), .Y(dp.rf._abc_6362_n3348) );
	NAND2X1 NAND2X1_1559 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n2975), .Y(dp.rf._abc_6362_n3070) );
	NAND2X1 NAND2X1_1560 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_17_<31>), .B(dp.rf._abc_6362_n2977), .Y(dp.rf._abc_6362_n3071_1) );
	NAND2X1 NAND2X1_1561 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3070), .B(dp.rf._abc_6362_n3071_1), .Y(dp.rf._abc_6362_n3349) );
	NAND2X1 NAND2X1_1562 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2172), .B(dp.rf._abc_6362_n2273), .Y(dp.rf._abc_6362_n3073_1) );
	NOR2X1 NOR2X1_200 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n3073_1), .Y(dp.rf._abc_6362_n3074) );
	NAND2X1 NAND2X1_1563 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3075_1) );
	INVX8 INVX8_14 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3076) );
	NAND2X1 NAND2X1_1564 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<0>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3077_1) );
	NAND2X1 NAND2X1_1565 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3075_1), .B(dp.rf._abc_6362_n3077_1), .Y(dp.rf._abc_6362_n3350) );
	NAND2X1 NAND2X1_1566 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3079_1) );
	NAND2X1 NAND2X1_1567 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<1>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3080) );
	NAND2X1 NAND2X1_1568 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3079_1), .B(dp.rf._abc_6362_n3080), .Y(dp.rf._abc_6362_n3351) );
	NAND2X1 NAND2X1_1569 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3082) );
	NAND2X1 NAND2X1_1570 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<2>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3083_1) );
	NAND2X1 NAND2X1_1571 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3082), .B(dp.rf._abc_6362_n3083_1), .Y(dp.rf._abc_6362_n3352) );
	NAND2X1 NAND2X1_1572 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3085_1) );
	NAND2X1 NAND2X1_1573 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<3>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3086) );
	NAND2X1 NAND2X1_1574 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3085_1), .B(dp.rf._abc_6362_n3086), .Y(dp.rf._abc_6362_n3353) );
	NAND2X1 NAND2X1_1575 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3088) );
	NAND2X1 NAND2X1_1576 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<4>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3089_1) );
	NAND2X1 NAND2X1_1577 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3088), .B(dp.rf._abc_6362_n3089_1), .Y(dp.rf._abc_6362_n3354) );
	NAND2X1 NAND2X1_1578 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3091_1) );
	NAND2X1 NAND2X1_1579 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<5>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3092) );
	NAND2X1 NAND2X1_1580 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3091_1), .B(dp.rf._abc_6362_n3092), .Y(dp.rf._abc_6362_n3355) );
	NAND2X1 NAND2X1_1581 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3094_1) );
	NAND2X1 NAND2X1_1582 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<6>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3095_1) );
	NAND2X1 NAND2X1_1583 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3094_1), .B(dp.rf._abc_6362_n3095_1), .Y(dp.rf._abc_6362_n3356) );
	NAND2X1 NAND2X1_1584 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3097_1) );
	NAND2X1 NAND2X1_1585 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<7>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3098_1) );
	NAND2X1 NAND2X1_1586 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3097_1), .B(dp.rf._abc_6362_n3098_1), .Y(dp.rf._abc_6362_n3357) );
	NAND2X1 NAND2X1_1587 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3100_1) );
	NAND2X1 NAND2X1_1588 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<8>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3101_1) );
	NAND2X1 NAND2X1_1589 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3100_1), .B(dp.rf._abc_6362_n3101_1), .Y(dp.rf._abc_6362_n3358) );
	NAND2X1 NAND2X1_1590 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3103_1) );
	NAND2X1 NAND2X1_1591 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<9>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3104_1) );
	NAND2X1 NAND2X1_1592 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3103_1), .B(dp.rf._abc_6362_n3104_1), .Y(dp.rf._abc_6362_n3359) );
	NAND2X1 NAND2X1_1593 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3106_1) );
	NAND2X1 NAND2X1_1594 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<10>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3107_1) );
	NAND2X1 NAND2X1_1595 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3106_1), .B(dp.rf._abc_6362_n3107_1), .Y(dp.rf._abc_6362_n3360) );
	NAND2X1 NAND2X1_1596 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3109_1) );
	NAND2X1 NAND2X1_1597 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<11>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3110_1) );
	NAND2X1 NAND2X1_1598 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3109_1), .B(dp.rf._abc_6362_n3110_1), .Y(dp.rf._abc_6362_n3361) );
	NAND2X1 NAND2X1_1599 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3112_1) );
	NAND2X1 NAND2X1_1600 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<12>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3113_1) );
	NAND2X1 NAND2X1_1601 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3112_1), .B(dp.rf._abc_6362_n3113_1), .Y(dp.rf._abc_6362_n3362) );
	NAND2X1 NAND2X1_1602 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3115_1) );
	NAND2X1 NAND2X1_1603 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<13>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3116_1) );
	NAND2X1 NAND2X1_1604 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3115_1), .B(dp.rf._abc_6362_n3116_1), .Y(dp.rf._abc_6362_n3363) );
	NAND2X1 NAND2X1_1605 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3118_1) );
	NAND2X1 NAND2X1_1606 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<14>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3119_1) );
	NAND2X1 NAND2X1_1607 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3118_1), .B(dp.rf._abc_6362_n3119_1), .Y(dp.rf._abc_6362_n3364) );
	NAND2X1 NAND2X1_1608 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3121_1) );
	NAND2X1 NAND2X1_1609 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<15>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3122_1) );
	NAND2X1 NAND2X1_1610 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3121_1), .B(dp.rf._abc_6362_n3122_1), .Y(dp.rf._abc_6362_n3365) );
	NAND2X1 NAND2X1_1611 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3124_1) );
	NAND2X1 NAND2X1_1612 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<16>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3125_1) );
	NAND2X1 NAND2X1_1613 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3124_1), .B(dp.rf._abc_6362_n3125_1), .Y(dp.rf._abc_6362_n3366) );
	NAND2X1 NAND2X1_1614 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3127_1) );
	NAND2X1 NAND2X1_1615 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<17>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3128_1) );
	NAND2X1 NAND2X1_1616 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3127_1), .B(dp.rf._abc_6362_n3128_1), .Y(dp.rf._abc_6362_n3367) );
	NAND2X1 NAND2X1_1617 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3130_1) );
	NAND2X1 NAND2X1_1618 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<18>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3131_1) );
	NAND2X1 NAND2X1_1619 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3130_1), .B(dp.rf._abc_6362_n3131_1), .Y(dp.rf._abc_6362_n3368) );
	NAND2X1 NAND2X1_1620 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3133_1) );
	NAND2X1 NAND2X1_1621 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<19>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3134_1) );
	NAND2X1 NAND2X1_1622 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3133_1), .B(dp.rf._abc_6362_n3134_1), .Y(dp.rf._abc_6362_n3369) );
	NAND2X1 NAND2X1_1623 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3136_1) );
	NAND2X1 NAND2X1_1624 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<20>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3137_1) );
	NAND2X1 NAND2X1_1625 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3136_1), .B(dp.rf._abc_6362_n3137_1), .Y(dp.rf._abc_6362_n3370) );
	NAND2X1 NAND2X1_1626 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3139_1) );
	NAND2X1 NAND2X1_1627 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<21>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3140_1) );
	NAND2X1 NAND2X1_1628 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3139_1), .B(dp.rf._abc_6362_n3140_1), .Y(dp.rf._abc_6362_n3371) );
	NAND2X1 NAND2X1_1629 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3142_1) );
	NAND2X1 NAND2X1_1630 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<22>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3143_1) );
	NAND2X1 NAND2X1_1631 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3142_1), .B(dp.rf._abc_6362_n3143_1), .Y(dp.rf._abc_6362_n3372) );
	NAND2X1 NAND2X1_1632 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3145_1) );
	NAND2X1 NAND2X1_1633 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<23>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3146_1) );
	NAND2X1 NAND2X1_1634 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3145_1), .B(dp.rf._abc_6362_n3146_1), .Y(dp.rf._abc_6362_n3373) );
	NAND2X1 NAND2X1_1635 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3148_1) );
	NAND2X1 NAND2X1_1636 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<24>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3149_1) );
	NAND2X1 NAND2X1_1637 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3148_1), .B(dp.rf._abc_6362_n3149_1), .Y(dp.rf._abc_6362_n3374) );
	NAND2X1 NAND2X1_1638 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3151_1) );
	NAND2X1 NAND2X1_1639 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<25>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3152_1) );
	NAND2X1 NAND2X1_1640 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3151_1), .B(dp.rf._abc_6362_n3152_1), .Y(dp.rf._abc_6362_n3375) );
	NAND2X1 NAND2X1_1641 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3154_1) );
	NAND2X1 NAND2X1_1642 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<26>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3155_1) );
	NAND2X1 NAND2X1_1643 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3154_1), .B(dp.rf._abc_6362_n3155_1), .Y(dp.rf._abc_6362_n3376) );
	NAND2X1 NAND2X1_1644 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3157_1) );
	NAND2X1 NAND2X1_1645 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<27>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3158_1) );
	NAND2X1 NAND2X1_1646 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3157_1), .B(dp.rf._abc_6362_n3158_1), .Y(dp.rf._abc_6362_n3377) );
	NAND2X1 NAND2X1_1647 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3160_1) );
	NAND2X1 NAND2X1_1648 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<28>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3161_1) );
	NAND2X1 NAND2X1_1649 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3160_1), .B(dp.rf._abc_6362_n3161_1), .Y(dp.rf._abc_6362_n3378) );
	NAND2X1 NAND2X1_1650 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3163_1) );
	NAND2X1 NAND2X1_1651 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<29>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3164_1) );
	NAND2X1 NAND2X1_1652 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3163_1), .B(dp.rf._abc_6362_n3164_1), .Y(dp.rf._abc_6362_n3379) );
	NAND2X1 NAND2X1_1653 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3166_1) );
	NAND2X1 NAND2X1_1654 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<30>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3167_1) );
	NAND2X1 NAND2X1_1655 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3166_1), .B(dp.rf._abc_6362_n3167_1), .Y(dp.rf._abc_6362_n3380) );
	NAND2X1 NAND2X1_1656 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n3074), .Y(dp.rf._abc_6362_n3169_1) );
	NAND2X1 NAND2X1_1657 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<31>), .B(dp.rf._abc_6362_n3076), .Y(dp.rf._abc_6362_n3170_1) );
	NAND2X1 NAND2X1_1658 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3169_1), .B(dp.rf._abc_6362_n3170_1), .Y(dp.rf._abc_6362_n3381) );
	NAND2X1 NAND2X1_1659 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2172), .B(dp.rf._abc_6362_n2376), .Y(dp.rf._abc_6362_n3172_1) );
	NOR2X1 NOR2X1_201 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n3172_1), .Y(dp.rf._abc_6362_n3173_1) );
	NAND2X1 NAND2X1_1660 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3174_1) );
	INVX8 INVX8_15 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3175_1) );
	NAND2X1 NAND2X1_1661 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<0>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3176_1) );
	NAND2X1 NAND2X1_1662 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3174_1), .B(dp.rf._abc_6362_n3176_1), .Y(dp.rf._abc_6362_n3382) );
	NAND2X1 NAND2X1_1663 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3178_1) );
	NAND2X1 NAND2X1_1664 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<1>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3179_1) );
	NAND2X1 NAND2X1_1665 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3178_1), .B(dp.rf._abc_6362_n3179_1), .Y(dp.rf._abc_6362_n3383) );
	NAND2X1 NAND2X1_1666 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3181_1) );
	NAND2X1 NAND2X1_1667 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<2>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3182_1) );
	NAND2X1 NAND2X1_1668 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3181_1), .B(dp.rf._abc_6362_n3182_1), .Y(dp.rf._abc_6362_n3384) );
	NAND2X1 NAND2X1_1669 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3184_1) );
	NAND2X1 NAND2X1_1670 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<3>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3185_1) );
	NAND2X1 NAND2X1_1671 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3184_1), .B(dp.rf._abc_6362_n3185_1), .Y(dp.rf._abc_6362_n3385) );
	NAND2X1 NAND2X1_1672 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3187_1) );
	NAND2X1 NAND2X1_1673 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<4>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3188_1) );
	NAND2X1 NAND2X1_1674 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3187_1), .B(dp.rf._abc_6362_n3188_1), .Y(dp.rf._abc_6362_n3386) );
	NAND2X1 NAND2X1_1675 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3190_1) );
	NAND2X1 NAND2X1_1676 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<5>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3191_1) );
	NAND2X1 NAND2X1_1677 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3190_1), .B(dp.rf._abc_6362_n3191_1), .Y(dp.rf._abc_6362_n3387) );
	NAND2X1 NAND2X1_1678 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3193_1) );
	NAND2X1 NAND2X1_1679 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<6>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3194_1) );
	NAND2X1 NAND2X1_1680 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3193_1), .B(dp.rf._abc_6362_n3194_1), .Y(dp.rf._abc_6362_n3388) );
	NAND2X1 NAND2X1_1681 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3196_1) );
	NAND2X1 NAND2X1_1682 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<7>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3197_1) );
	NAND2X1 NAND2X1_1683 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3196_1), .B(dp.rf._abc_6362_n3197_1), .Y(dp.rf._abc_6362_n3389) );
	NAND2X1 NAND2X1_1684 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3199_1) );
	NAND2X1 NAND2X1_1685 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<8>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3200_1) );
	NAND2X1 NAND2X1_1686 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3199_1), .B(dp.rf._abc_6362_n3200_1), .Y(dp.rf._abc_6362_n3390) );
	NAND2X1 NAND2X1_1687 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3202_1) );
	NAND2X1 NAND2X1_1688 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<9>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3203_1) );
	NAND2X1 NAND2X1_1689 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3202_1), .B(dp.rf._abc_6362_n3203_1), .Y(dp.rf._abc_6362_n3391) );
	NAND2X1 NAND2X1_1690 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3205_1) );
	NAND2X1 NAND2X1_1691 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<10>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3206_1) );
	NAND2X1 NAND2X1_1692 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3205_1), .B(dp.rf._abc_6362_n3206_1), .Y(dp.rf._abc_6362_n3392) );
	NAND2X1 NAND2X1_1693 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3208_1) );
	NAND2X1 NAND2X1_1694 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<11>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3209_1) );
	NAND2X1 NAND2X1_1695 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3208_1), .B(dp.rf._abc_6362_n3209_1), .Y(dp.rf._abc_6362_n3393) );
	NAND2X1 NAND2X1_1696 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3211_1) );
	NAND2X1 NAND2X1_1697 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<12>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3212_1) );
	NAND2X1 NAND2X1_1698 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3211_1), .B(dp.rf._abc_6362_n3212_1), .Y(dp.rf._abc_6362_n3394) );
	NAND2X1 NAND2X1_1699 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3214_1) );
	NAND2X1 NAND2X1_1700 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<13>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3215_1) );
	NAND2X1 NAND2X1_1701 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3214_1), .B(dp.rf._abc_6362_n3215_1), .Y(dp.rf._abc_6362_n3395) );
	NAND2X1 NAND2X1_1702 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3217_1) );
	NAND2X1 NAND2X1_1703 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<14>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3218_1) );
	NAND2X1 NAND2X1_1704 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3217_1), .B(dp.rf._abc_6362_n3218_1), .Y(dp.rf._abc_6362_n3396) );
	NAND2X1 NAND2X1_1705 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3220_1) );
	NAND2X1 NAND2X1_1706 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<15>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3221_1) );
	NAND2X1 NAND2X1_1707 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3220_1), .B(dp.rf._abc_6362_n3221_1), .Y(dp.rf._abc_6362_n3397) );
	NAND2X1 NAND2X1_1708 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3223_1) );
	NAND2X1 NAND2X1_1709 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<16>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3224_1) );
	NAND2X1 NAND2X1_1710 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3223_1), .B(dp.rf._abc_6362_n3224_1), .Y(dp.rf._abc_6362_n3398) );
	NAND2X1 NAND2X1_1711 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3226_1) );
	NAND2X1 NAND2X1_1712 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<17>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3227_1) );
	NAND2X1 NAND2X1_1713 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3226_1), .B(dp.rf._abc_6362_n3227_1), .Y(dp.rf._abc_6362_n3399) );
	NAND2X1 NAND2X1_1714 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3229_1) );
	NAND2X1 NAND2X1_1715 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<18>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3230_1) );
	NAND2X1 NAND2X1_1716 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3229_1), .B(dp.rf._abc_6362_n3230_1), .Y(dp.rf._abc_6362_n3400) );
	NAND2X1 NAND2X1_1717 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3232_1) );
	NAND2X1 NAND2X1_1718 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<19>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3233_1) );
	NAND2X1 NAND2X1_1719 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3232_1), .B(dp.rf._abc_6362_n3233_1), .Y(dp.rf._abc_6362_n3401) );
	NAND2X1 NAND2X1_1720 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3235_1) );
	NAND2X1 NAND2X1_1721 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<20>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3236_1) );
	NAND2X1 NAND2X1_1722 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3235_1), .B(dp.rf._abc_6362_n3236_1), .Y(dp.rf._abc_6362_n3402) );
	NAND2X1 NAND2X1_1723 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3238_1) );
	NAND2X1 NAND2X1_1724 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<21>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3239_1) );
	NAND2X1 NAND2X1_1725 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3238_1), .B(dp.rf._abc_6362_n3239_1), .Y(dp.rf._abc_6362_n3403) );
	NAND2X1 NAND2X1_1726 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3241_1) );
	NAND2X1 NAND2X1_1727 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<22>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3242_1) );
	NAND2X1 NAND2X1_1728 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3241_1), .B(dp.rf._abc_6362_n3242_1), .Y(dp.rf._abc_6362_n3404) );
	NAND2X1 NAND2X1_1729 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3244_1) );
	NAND2X1 NAND2X1_1730 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<23>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3245_1) );
	NAND2X1 NAND2X1_1731 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3244_1), .B(dp.rf._abc_6362_n3245_1), .Y(dp.rf._abc_6362_n3405) );
	NAND2X1 NAND2X1_1732 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3247_1) );
	NAND2X1 NAND2X1_1733 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<24>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3248_1) );
	NAND2X1 NAND2X1_1734 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3247_1), .B(dp.rf._abc_6362_n3248_1), .Y(dp.rf._abc_6362_n3406) );
	NAND2X1 NAND2X1_1735 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3250_1) );
	NAND2X1 NAND2X1_1736 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<25>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3251_1) );
	NAND2X1 NAND2X1_1737 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3250_1), .B(dp.rf._abc_6362_n3251_1), .Y(dp.rf._abc_6362_n3407) );
	NAND2X1 NAND2X1_1738 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3253_1) );
	NAND2X1 NAND2X1_1739 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<26>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3254_1) );
	NAND2X1 NAND2X1_1740 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3253_1), .B(dp.rf._abc_6362_n3254_1), .Y(dp.rf._abc_6362_n3408) );
	NAND2X1 NAND2X1_1741 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3256_1) );
	NAND2X1 NAND2X1_1742 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<27>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3257_1) );
	NAND2X1 NAND2X1_1743 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3256_1), .B(dp.rf._abc_6362_n3257_1), .Y(dp.rf._abc_6362_n3409) );
	NAND2X1 NAND2X1_1744 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3259_1) );
	NAND2X1 NAND2X1_1745 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<28>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3260_1) );
	NAND2X1 NAND2X1_1746 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3259_1), .B(dp.rf._abc_6362_n3260_1), .Y(dp.rf._abc_6362_n3410) );
	NAND2X1 NAND2X1_1747 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3262_1) );
	NAND2X1 NAND2X1_1748 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<29>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3263_1) );
	NAND2X1 NAND2X1_1749 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3262_1), .B(dp.rf._abc_6362_n3263_1), .Y(dp.rf._abc_6362_n3411) );
	NAND2X1 NAND2X1_1750 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3265_1) );
	NAND2X1 NAND2X1_1751 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<30>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3266_1) );
	NAND2X1 NAND2X1_1752 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3265_1), .B(dp.rf._abc_6362_n3266_1), .Y(dp.rf._abc_6362_n3412) );
	NAND2X1 NAND2X1_1753 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n3173_1), .Y(dp.rf._abc_6362_n3268_1) );
	NAND2X1 NAND2X1_1754 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_19_<31>), .B(dp.rf._abc_6362_n3175_1), .Y(dp.rf._abc_6362_n3269_1) );
	NAND2X1 NAND2X1_1755 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3268_1), .B(dp.rf._abc_6362_n3269_1), .Y(dp.rf._abc_6362_n3413) );
	NOR2X1 NOR2X1_202 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n2974), .Y(dp.rf._abc_6362_n3271_1) );
	NAND2X1 NAND2X1_1756 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3272_1) );
	INVX8 INVX8_16 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3273_1) );
	NAND2X1 NAND2X1_1757 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<0>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3274_1) );
	NAND2X1 NAND2X1_1758 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3272_1), .B(dp.rf._abc_6362_n3274_1), .Y(dp.rf._abc_6362_n3414) );
	NAND2X1 NAND2X1_1759 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3276_1) );
	NAND2X1 NAND2X1_1760 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<1>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3277_1) );
	NAND2X1 NAND2X1_1761 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3276_1), .B(dp.rf._abc_6362_n3277_1), .Y(dp.rf._abc_6362_n3415) );
	NAND2X1 NAND2X1_1762 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3279_1) );
	NAND2X1 NAND2X1_1763 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<2>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3280_1) );
	NAND2X1 NAND2X1_1764 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3279_1), .B(dp.rf._abc_6362_n3280_1), .Y(dp.rf._abc_6362_n3416) );
	NAND2X1 NAND2X1_1765 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3282_1) );
	NAND2X1 NAND2X1_1766 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<3>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3283_1) );
	NAND2X1 NAND2X1_1767 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3282_1), .B(dp.rf._abc_6362_n3283_1), .Y(dp.rf._abc_6362_n3417) );
	NAND2X1 NAND2X1_1768 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3285_1) );
	NAND2X1 NAND2X1_1769 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<4>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3286_1) );
	NAND2X1 NAND2X1_1770 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3285_1), .B(dp.rf._abc_6362_n3286_1), .Y(dp.rf._abc_6362_n3418) );
	NAND2X1 NAND2X1_1771 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3288_1) );
	NAND2X1 NAND2X1_1772 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<5>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3289_1) );
	NAND2X1 NAND2X1_1773 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3288_1), .B(dp.rf._abc_6362_n3289_1), .Y(dp.rf._abc_6362_n3419) );
	NAND2X1 NAND2X1_1774 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3291_1) );
	NAND2X1 NAND2X1_1775 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<6>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3292_1) );
	NAND2X1 NAND2X1_1776 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3291_1), .B(dp.rf._abc_6362_n3292_1), .Y(dp.rf._abc_6362_n3420) );
	NAND2X1 NAND2X1_1777 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3294_1) );
	NAND2X1 NAND2X1_1778 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<7>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3295_1) );
	NAND2X1 NAND2X1_1779 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3294_1), .B(dp.rf._abc_6362_n3295_1), .Y(dp.rf._abc_6362_n3421) );
	NAND2X1 NAND2X1_1780 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3297_1) );
	NAND2X1 NAND2X1_1781 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<8>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3298_1) );
	NAND2X1 NAND2X1_1782 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3297_1), .B(dp.rf._abc_6362_n3298_1), .Y(dp.rf._abc_6362_n3422) );
	NAND2X1 NAND2X1_1783 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3300_1) );
	NAND2X1 NAND2X1_1784 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<9>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3301_1) );
	NAND2X1 NAND2X1_1785 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3300_1), .B(dp.rf._abc_6362_n3301_1), .Y(dp.rf._abc_6362_n3423) );
	NAND2X1 NAND2X1_1786 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3303_1) );
	NAND2X1 NAND2X1_1787 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<10>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3304_1) );
	NAND2X1 NAND2X1_1788 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3303_1), .B(dp.rf._abc_6362_n3304_1), .Y(dp.rf._abc_6362_n3424) );
	NAND2X1 NAND2X1_1789 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3306_1) );
	NAND2X1 NAND2X1_1790 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<11>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3307_1) );
	NAND2X1 NAND2X1_1791 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3306_1), .B(dp.rf._abc_6362_n3307_1), .Y(dp.rf._abc_6362_n3425) );
	NAND2X1 NAND2X1_1792 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3309_1) );
	NAND2X1 NAND2X1_1793 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<12>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3310_1) );
	NAND2X1 NAND2X1_1794 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3309_1), .B(dp.rf._abc_6362_n3310_1), .Y(dp.rf._abc_6362_n3426) );
	NAND2X1 NAND2X1_1795 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3312_1) );
	NAND2X1 NAND2X1_1796 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<13>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3313_1) );
	NAND2X1 NAND2X1_1797 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3312_1), .B(dp.rf._abc_6362_n3313_1), .Y(dp.rf._abc_6362_n3427) );
	NAND2X1 NAND2X1_1798 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3315_1) );
	NAND2X1 NAND2X1_1799 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<14>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3316_1) );
	NAND2X1 NAND2X1_1800 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3315_1), .B(dp.rf._abc_6362_n3316_1), .Y(dp.rf._abc_6362_n3428) );
	NAND2X1 NAND2X1_1801 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3318_1) );
	NAND2X1 NAND2X1_1802 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<15>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3319_1) );
	NAND2X1 NAND2X1_1803 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3318_1), .B(dp.rf._abc_6362_n3319_1), .Y(dp.rf._abc_6362_n3429) );
	NAND2X1 NAND2X1_1804 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3321_1) );
	NAND2X1 NAND2X1_1805 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<16>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3322_1) );
	NAND2X1 NAND2X1_1806 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3321_1), .B(dp.rf._abc_6362_n3322_1), .Y(dp.rf._abc_6362_n3430) );
	NAND2X1 NAND2X1_1807 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3324_1) );
	NAND2X1 NAND2X1_1808 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<17>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3325_1) );
	NAND2X1 NAND2X1_1809 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3324_1), .B(dp.rf._abc_6362_n3325_1), .Y(dp.rf._abc_6362_n3431) );
	NAND2X1 NAND2X1_1810 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3327_1) );
	NAND2X1 NAND2X1_1811 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<18>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3328_1) );
	NAND2X1 NAND2X1_1812 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3327_1), .B(dp.rf._abc_6362_n3328_1), .Y(dp.rf._abc_6362_n3432) );
	NAND2X1 NAND2X1_1813 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3330_1) );
	NAND2X1 NAND2X1_1814 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<19>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3331_1) );
	NAND2X1 NAND2X1_1815 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3330_1), .B(dp.rf._abc_6362_n3331_1), .Y(dp.rf._abc_6362_n3433) );
	NAND2X1 NAND2X1_1816 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3333_1) );
	NAND2X1 NAND2X1_1817 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<20>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3334_1) );
	NAND2X1 NAND2X1_1818 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3333_1), .B(dp.rf._abc_6362_n3334_1), .Y(dp.rf._abc_6362_n3434) );
	NAND2X1 NAND2X1_1819 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3336_1) );
	NAND2X1 NAND2X1_1820 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<21>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3337_1) );
	NAND2X1 NAND2X1_1821 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3336_1), .B(dp.rf._abc_6362_n3337_1), .Y(dp.rf._abc_6362_n3435) );
	NAND2X1 NAND2X1_1822 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3339_1) );
	NAND2X1 NAND2X1_1823 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<22>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3340_1) );
	NAND2X1 NAND2X1_1824 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3339_1), .B(dp.rf._abc_6362_n3340_1), .Y(dp.rf._abc_6362_n3436) );
	NAND2X1 NAND2X1_1825 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3342_1) );
	NAND2X1 NAND2X1_1826 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<23>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3343_1) );
	NAND2X1 NAND2X1_1827 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3342_1), .B(dp.rf._abc_6362_n3343_1), .Y(dp.rf._abc_6362_n3437) );
	NAND2X1 NAND2X1_1828 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3345_1) );
	NAND2X1 NAND2X1_1829 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<24>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3346_1) );
	NAND2X1 NAND2X1_1830 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3345_1), .B(dp.rf._abc_6362_n3346_1), .Y(dp.rf._abc_6362_n3438) );
	NAND2X1 NAND2X1_1831 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3348_1) );
	NAND2X1 NAND2X1_1832 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<25>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3349_1) );
	NAND2X1 NAND2X1_1833 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3348_1), .B(dp.rf._abc_6362_n3349_1), .Y(dp.rf._abc_6362_n3439) );
	NAND2X1 NAND2X1_1834 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3351_1) );
	NAND2X1 NAND2X1_1835 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<26>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3352_1) );
	NAND2X1 NAND2X1_1836 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3351_1), .B(dp.rf._abc_6362_n3352_1), .Y(dp.rf._abc_6362_n3440) );
	NAND2X1 NAND2X1_1837 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3354_1) );
	NAND2X1 NAND2X1_1838 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<27>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3355_1) );
	NAND2X1 NAND2X1_1839 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3354_1), .B(dp.rf._abc_6362_n3355_1), .Y(dp.rf._abc_6362_n3441) );
	NAND2X1 NAND2X1_1840 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3357_1) );
	NAND2X1 NAND2X1_1841 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<28>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3358_1) );
	NAND2X1 NAND2X1_1842 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3357_1), .B(dp.rf._abc_6362_n3358_1), .Y(dp.rf._abc_6362_n3442) );
	NAND2X1 NAND2X1_1843 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3360_1) );
	NAND2X1 NAND2X1_1844 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<29>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3361_1) );
	NAND2X1 NAND2X1_1845 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3360_1), .B(dp.rf._abc_6362_n3361_1), .Y(dp.rf._abc_6362_n3443) );
	NAND2X1 NAND2X1_1846 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3363_1) );
	NAND2X1 NAND2X1_1847 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<30>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3364_1) );
	NAND2X1 NAND2X1_1848 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3363_1), .B(dp.rf._abc_6362_n3364_1), .Y(dp.rf._abc_6362_n3444) );
	NAND2X1 NAND2X1_1849 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n3271_1), .Y(dp.rf._abc_6362_n3366_1) );
	NAND2X1 NAND2X1_1850 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<31>), .B(dp.rf._abc_6362_n3273_1), .Y(dp.rf._abc_6362_n3367_1) );
	NAND2X1 NAND2X1_1851 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3366_1), .B(dp.rf._abc_6362_n3367_1), .Y(dp.rf._abc_6362_n3445) );
	NAND2X1 NAND2X1_1852 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2170), .B(dp.rf._abc_6362_n2169), .Y(dp.rf._abc_6362_n3369_1) );
	INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3369_1), .Y(dp.rf._abc_6362_n3370_1) );
	NAND2X1 NAND2X1_1853 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2167), .B(dp.rf._abc_6362_n3370_1), .Y(dp.rf._abc_6362_n3371_1) );
	NOR2X1 NOR2X1_203 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n3371_1), .Y(dp.rf._abc_6362_n3372_1) );
	NAND2X1 NAND2X1_1854 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3373_1) );
	INVX8 INVX8_17 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3374_1) );
	NAND2X1 NAND2X1_1855 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<0>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3375_1) );
	NAND2X1 NAND2X1_1856 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3373_1), .B(dp.rf._abc_6362_n3375_1), .Y(dp.rf._abc_6362_n3446) );
	NAND2X1 NAND2X1_1857 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3377_1) );
	NAND2X1 NAND2X1_1858 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<1>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3378_1) );
	NAND2X1 NAND2X1_1859 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3377_1), .B(dp.rf._abc_6362_n3378_1), .Y(dp.rf._abc_6362_n3447) );
	NAND2X1 NAND2X1_1860 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3380_1) );
	NAND2X1 NAND2X1_1861 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<2>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3381_1) );
	NAND2X1 NAND2X1_1862 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3380_1), .B(dp.rf._abc_6362_n3381_1), .Y(dp.rf._abc_6362_n3448) );
	NAND2X1 NAND2X1_1863 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3383_1) );
	NAND2X1 NAND2X1_1864 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<3>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3384_1) );
	NAND2X1 NAND2X1_1865 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3383_1), .B(dp.rf._abc_6362_n3384_1), .Y(dp.rf._abc_6362_n3449) );
	NAND2X1 NAND2X1_1866 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3386_1) );
	NAND2X1 NAND2X1_1867 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<4>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3387_1) );
	NAND2X1 NAND2X1_1868 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3386_1), .B(dp.rf._abc_6362_n3387_1), .Y(dp.rf._abc_6362_n3450) );
	NAND2X1 NAND2X1_1869 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3389_1) );
	NAND2X1 NAND2X1_1870 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<5>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3390_1) );
	NAND2X1 NAND2X1_1871 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3389_1), .B(dp.rf._abc_6362_n3390_1), .Y(dp.rf._abc_6362_n3451) );
	NAND2X1 NAND2X1_1872 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3392_1) );
	NAND2X1 NAND2X1_1873 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<6>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3393_1) );
	NAND2X1 NAND2X1_1874 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3392_1), .B(dp.rf._abc_6362_n3393_1), .Y(dp.rf._abc_6362_n3452) );
	NAND2X1 NAND2X1_1875 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3395_1) );
	NAND2X1 NAND2X1_1876 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<7>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3396_1) );
	NAND2X1 NAND2X1_1877 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3395_1), .B(dp.rf._abc_6362_n3396_1), .Y(dp.rf._abc_6362_n3453) );
	NAND2X1 NAND2X1_1878 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3398_1) );
	NAND2X1 NAND2X1_1879 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<8>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3399_1) );
	NAND2X1 NAND2X1_1880 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3398_1), .B(dp.rf._abc_6362_n3399_1), .Y(dp.rf._abc_6362_n3454) );
	NAND2X1 NAND2X1_1881 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3401_1) );
	NAND2X1 NAND2X1_1882 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<9>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3402_1) );
	NAND2X1 NAND2X1_1883 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3401_1), .B(dp.rf._abc_6362_n3402_1), .Y(dp.rf._abc_6362_n3455) );
	NAND2X1 NAND2X1_1884 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3404_1) );
	NAND2X1 NAND2X1_1885 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<10>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3405_1) );
	NAND2X1 NAND2X1_1886 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3404_1), .B(dp.rf._abc_6362_n3405_1), .Y(dp.rf._abc_6362_n3456) );
	NAND2X1 NAND2X1_1887 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3407_1) );
	NAND2X1 NAND2X1_1888 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<11>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3408_1) );
	NAND2X1 NAND2X1_1889 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3407_1), .B(dp.rf._abc_6362_n3408_1), .Y(dp.rf._abc_6362_n3457) );
	NAND2X1 NAND2X1_1890 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3410_1) );
	NAND2X1 NAND2X1_1891 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<12>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3411_1) );
	NAND2X1 NAND2X1_1892 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3410_1), .B(dp.rf._abc_6362_n3411_1), .Y(dp.rf._abc_6362_n3458) );
	NAND2X1 NAND2X1_1893 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3413_1) );
	NAND2X1 NAND2X1_1894 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<13>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3414_1) );
	NAND2X1 NAND2X1_1895 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3413_1), .B(dp.rf._abc_6362_n3414_1), .Y(dp.rf._abc_6362_n3459) );
	NAND2X1 NAND2X1_1896 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3416_1) );
	NAND2X1 NAND2X1_1897 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<14>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3417_1) );
	NAND2X1 NAND2X1_1898 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3416_1), .B(dp.rf._abc_6362_n3417_1), .Y(dp.rf._abc_6362_n3460) );
	NAND2X1 NAND2X1_1899 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3419_1) );
	NAND2X1 NAND2X1_1900 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<15>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3420_1) );
	NAND2X1 NAND2X1_1901 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3419_1), .B(dp.rf._abc_6362_n3420_1), .Y(dp.rf._abc_6362_n3461) );
	NAND2X1 NAND2X1_1902 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3422_1) );
	NAND2X1 NAND2X1_1903 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<16>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3423_1) );
	NAND2X1 NAND2X1_1904 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3422_1), .B(dp.rf._abc_6362_n3423_1), .Y(dp.rf._abc_6362_n3462) );
	NAND2X1 NAND2X1_1905 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3425_1) );
	NAND2X1 NAND2X1_1906 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<17>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3426_1) );
	NAND2X1 NAND2X1_1907 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3425_1), .B(dp.rf._abc_6362_n3426_1), .Y(dp.rf._abc_6362_n3463) );
	NAND2X1 NAND2X1_1908 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3428_1) );
	NAND2X1 NAND2X1_1909 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<18>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3429_1) );
	NAND2X1 NAND2X1_1910 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3428_1), .B(dp.rf._abc_6362_n3429_1), .Y(dp.rf._abc_6362_n3464) );
	NAND2X1 NAND2X1_1911 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3431_1) );
	NAND2X1 NAND2X1_1912 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<19>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3432_1) );
	NAND2X1 NAND2X1_1913 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3431_1), .B(dp.rf._abc_6362_n3432_1), .Y(dp.rf._abc_6362_n3465) );
	NAND2X1 NAND2X1_1914 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3434_1) );
	NAND2X1 NAND2X1_1915 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<20>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3435_1) );
	NAND2X1 NAND2X1_1916 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3434_1), .B(dp.rf._abc_6362_n3435_1), .Y(dp.rf._abc_6362_n3466) );
	NAND2X1 NAND2X1_1917 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3437_1) );
	NAND2X1 NAND2X1_1918 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<21>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3438_1) );
	NAND2X1 NAND2X1_1919 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3437_1), .B(dp.rf._abc_6362_n3438_1), .Y(dp.rf._abc_6362_n3467) );
	NAND2X1 NAND2X1_1920 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3440_1) );
	NAND2X1 NAND2X1_1921 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<22>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3441_1) );
	NAND2X1 NAND2X1_1922 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3440_1), .B(dp.rf._abc_6362_n3441_1), .Y(dp.rf._abc_6362_n3468) );
	NAND2X1 NAND2X1_1923 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3443_1) );
	NAND2X1 NAND2X1_1924 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<23>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3444_1) );
	NAND2X1 NAND2X1_1925 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3443_1), .B(dp.rf._abc_6362_n3444_1), .Y(dp.rf._abc_6362_n3469) );
	NAND2X1 NAND2X1_1926 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3446_1) );
	NAND2X1 NAND2X1_1927 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<24>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3447_1) );
	NAND2X1 NAND2X1_1928 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3446_1), .B(dp.rf._abc_6362_n3447_1), .Y(dp.rf._abc_6362_n3470) );
	NAND2X1 NAND2X1_1929 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3449_1) );
	NAND2X1 NAND2X1_1930 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<25>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3450_1) );
	NAND2X1 NAND2X1_1931 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3449_1), .B(dp.rf._abc_6362_n3450_1), .Y(dp.rf._abc_6362_n3471) );
	NAND2X1 NAND2X1_1932 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3452_1) );
	NAND2X1 NAND2X1_1933 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<26>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3453_1) );
	NAND2X1 NAND2X1_1934 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3452_1), .B(dp.rf._abc_6362_n3453_1), .Y(dp.rf._abc_6362_n3472) );
	NAND2X1 NAND2X1_1935 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3455_1) );
	NAND2X1 NAND2X1_1936 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<27>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3456_1) );
	NAND2X1 NAND2X1_1937 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3455_1), .B(dp.rf._abc_6362_n3456_1), .Y(dp.rf._abc_6362_n3473) );
	NAND2X1 NAND2X1_1938 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3458_1) );
	NAND2X1 NAND2X1_1939 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<28>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3459_1) );
	NAND2X1 NAND2X1_1940 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3458_1), .B(dp.rf._abc_6362_n3459_1), .Y(dp.rf._abc_6362_n3474) );
	NAND2X1 NAND2X1_1941 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3461_1) );
	NAND2X1 NAND2X1_1942 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<29>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3462_1) );
	NAND2X1 NAND2X1_1943 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3461_1), .B(dp.rf._abc_6362_n3462_1), .Y(dp.rf._abc_6362_n3475) );
	NAND2X1 NAND2X1_1944 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3464_1) );
	NAND2X1 NAND2X1_1945 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<30>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3465_1) );
	NAND2X1 NAND2X1_1946 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3464_1), .B(dp.rf._abc_6362_n3465_1), .Y(dp.rf._abc_6362_n3476) );
	NAND2X1 NAND2X1_1947 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n3372_1), .Y(dp.rf._abc_6362_n3467_1) );
	NAND2X1 NAND2X1_1948 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<31>), .B(dp.rf._abc_6362_n3374_1), .Y(dp.rf._abc_6362_n3468_1) );
	NAND2X1 NAND2X1_1949 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3467_1), .B(dp.rf._abc_6362_n3468_1), .Y(dp.rf._abc_6362_n3477) );
	NAND2X1 NAND2X1_1950 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3370_1), .B(dp.rf._abc_6362_n2576), .Y(dp.rf._abc_6362_n3470_1) );
	NOR2X1 NOR2X1_204 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n3470_1), .Y(dp.rf._abc_6362_n3471_1) );
	NAND2X1 NAND2X1_1951 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3472_1) );
	INVX8 INVX8_18 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3473_1) );
	NAND2X1 NAND2X1_1952 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<0>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3474_1) );
	NAND2X1 NAND2X1_1953 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3472_1), .B(dp.rf._abc_6362_n3474_1), .Y(dp.rf._abc_6362_n3478) );
	NAND2X1 NAND2X1_1954 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3476_1) );
	NAND2X1 NAND2X1_1955 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<1>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3477_1) );
	NAND2X1 NAND2X1_1956 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3476_1), .B(dp.rf._abc_6362_n3477_1), .Y(dp.rf._abc_6362_n3479) );
	NAND2X1 NAND2X1_1957 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3479_1) );
	NAND2X1 NAND2X1_1958 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<2>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3480_1) );
	NAND2X1 NAND2X1_1959 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3479_1), .B(dp.rf._abc_6362_n3480_1), .Y(dp.rf._abc_6362_n3480) );
	NAND2X1 NAND2X1_1960 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3482_1) );
	NAND2X1 NAND2X1_1961 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<3>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3483_1) );
	NAND2X1 NAND2X1_1962 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3482_1), .B(dp.rf._abc_6362_n3483_1), .Y(dp.rf._abc_6362_n3481) );
	NAND2X1 NAND2X1_1963 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3485_1) );
	NAND2X1 NAND2X1_1964 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<4>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3486_1) );
	NAND2X1 NAND2X1_1965 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3485_1), .B(dp.rf._abc_6362_n3486_1), .Y(dp.rf._abc_6362_n3482) );
	NAND2X1 NAND2X1_1966 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3488_1) );
	NAND2X1 NAND2X1_1967 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<5>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3489_1) );
	NAND2X1 NAND2X1_1968 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3488_1), .B(dp.rf._abc_6362_n3489_1), .Y(dp.rf._abc_6362_n3483) );
	NAND2X1 NAND2X1_1969 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3491_1) );
	NAND2X1 NAND2X1_1970 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<6>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3492_1) );
	NAND2X1 NAND2X1_1971 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3491_1), .B(dp.rf._abc_6362_n3492_1), .Y(dp.rf._abc_6362_n3484) );
	NAND2X1 NAND2X1_1972 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3494_1) );
	NAND2X1 NAND2X1_1973 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<7>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3495_1) );
	NAND2X1 NAND2X1_1974 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3494_1), .B(dp.rf._abc_6362_n3495_1), .Y(dp.rf._abc_6362_n3485) );
	NAND2X1 NAND2X1_1975 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3497_1) );
	NAND2X1 NAND2X1_1976 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<8>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3498_1) );
	NAND2X1 NAND2X1_1977 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3497_1), .B(dp.rf._abc_6362_n3498_1), .Y(dp.rf._abc_6362_n3486) );
	NAND2X1 NAND2X1_1978 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3500_1) );
	NAND2X1 NAND2X1_1979 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<9>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3501_1) );
	NAND2X1 NAND2X1_1980 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3500_1), .B(dp.rf._abc_6362_n3501_1), .Y(dp.rf._abc_6362_n3487) );
	NAND2X1 NAND2X1_1981 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3503_1) );
	NAND2X1 NAND2X1_1982 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<10>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3504_1) );
	NAND2X1 NAND2X1_1983 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3503_1), .B(dp.rf._abc_6362_n3504_1), .Y(dp.rf._abc_6362_n3488) );
	NAND2X1 NAND2X1_1984 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3506_1) );
	NAND2X1 NAND2X1_1985 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<11>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3507_1) );
	NAND2X1 NAND2X1_1986 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3506_1), .B(dp.rf._abc_6362_n3507_1), .Y(dp.rf._abc_6362_n3489) );
	NAND2X1 NAND2X1_1987 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3509_1) );
	NAND2X1 NAND2X1_1988 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<12>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3510_1) );
	NAND2X1 NAND2X1_1989 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3509_1), .B(dp.rf._abc_6362_n3510_1), .Y(dp.rf._abc_6362_n3490) );
	NAND2X1 NAND2X1_1990 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3512_1) );
	NAND2X1 NAND2X1_1991 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<13>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3513_1) );
	NAND2X1 NAND2X1_1992 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3512_1), .B(dp.rf._abc_6362_n3513_1), .Y(dp.rf._abc_6362_n3491) );
	NAND2X1 NAND2X1_1993 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3515_1) );
	NAND2X1 NAND2X1_1994 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<14>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3516_1) );
	NAND2X1 NAND2X1_1995 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3515_1), .B(dp.rf._abc_6362_n3516_1), .Y(dp.rf._abc_6362_n3492) );
	NAND2X1 NAND2X1_1996 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3518_1) );
	NAND2X1 NAND2X1_1997 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<15>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3519_1) );
	NAND2X1 NAND2X1_1998 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3518_1), .B(dp.rf._abc_6362_n3519_1), .Y(dp.rf._abc_6362_n3493) );
	NAND2X1 NAND2X1_1999 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3521_1) );
	NAND2X1 NAND2X1_2000 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<16>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3522_1) );
	NAND2X1 NAND2X1_2001 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3521_1), .B(dp.rf._abc_6362_n3522_1), .Y(dp.rf._abc_6362_n3494) );
	NAND2X1 NAND2X1_2002 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3524_1) );
	NAND2X1 NAND2X1_2003 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<17>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3525_1) );
	NAND2X1 NAND2X1_2004 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3524_1), .B(dp.rf._abc_6362_n3525_1), .Y(dp.rf._abc_6362_n3495) );
	NAND2X1 NAND2X1_2005 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3527_1) );
	NAND2X1 NAND2X1_2006 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<18>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3528_1) );
	NAND2X1 NAND2X1_2007 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3527_1), .B(dp.rf._abc_6362_n3528_1), .Y(dp.rf._abc_6362_n3496) );
	NAND2X1 NAND2X1_2008 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3530_1) );
	NAND2X1 NAND2X1_2009 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<19>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3531_1) );
	NAND2X1 NAND2X1_2010 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3530_1), .B(dp.rf._abc_6362_n3531_1), .Y(dp.rf._abc_6362_n3497) );
	NAND2X1 NAND2X1_2011 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3533_1) );
	NAND2X1 NAND2X1_2012 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<20>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3534_1) );
	NAND2X1 NAND2X1_2013 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3533_1), .B(dp.rf._abc_6362_n3534_1), .Y(dp.rf._abc_6362_n3498) );
	NAND2X1 NAND2X1_2014 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3536_1) );
	NAND2X1 NAND2X1_2015 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<21>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3537_1) );
	NAND2X1 NAND2X1_2016 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3536_1), .B(dp.rf._abc_6362_n3537_1), .Y(dp.rf._abc_6362_n3499) );
	NAND2X1 NAND2X1_2017 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3539_1) );
	NAND2X1 NAND2X1_2018 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<22>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3540_1) );
	NAND2X1 NAND2X1_2019 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3539_1), .B(dp.rf._abc_6362_n3540_1), .Y(dp.rf._abc_6362_n3500) );
	NAND2X1 NAND2X1_2020 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3542_1) );
	NAND2X1 NAND2X1_2021 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<23>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3543_1) );
	NAND2X1 NAND2X1_2022 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3542_1), .B(dp.rf._abc_6362_n3543_1), .Y(dp.rf._abc_6362_n3501) );
	NAND2X1 NAND2X1_2023 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3545_1) );
	NAND2X1 NAND2X1_2024 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<24>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3546_1) );
	NAND2X1 NAND2X1_2025 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3545_1), .B(dp.rf._abc_6362_n3546_1), .Y(dp.rf._abc_6362_n3502) );
	NAND2X1 NAND2X1_2026 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3548_1) );
	NAND2X1 NAND2X1_2027 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<25>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3549_1) );
	NAND2X1 NAND2X1_2028 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3548_1), .B(dp.rf._abc_6362_n3549_1), .Y(dp.rf._abc_6362_n3503) );
	NAND2X1 NAND2X1_2029 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3551_1) );
	NAND2X1 NAND2X1_2030 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<26>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3552_1) );
	NAND2X1 NAND2X1_2031 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3551_1), .B(dp.rf._abc_6362_n3552_1), .Y(dp.rf._abc_6362_n3504) );
	NAND2X1 NAND2X1_2032 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3554_1) );
	NAND2X1 NAND2X1_2033 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<27>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3555_1) );
	NAND2X1 NAND2X1_2034 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3554_1), .B(dp.rf._abc_6362_n3555_1), .Y(dp.rf._abc_6362_n3505) );
	NAND2X1 NAND2X1_2035 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3557_1) );
	NAND2X1 NAND2X1_2036 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<28>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3558_1) );
	NAND2X1 NAND2X1_2037 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3557_1), .B(dp.rf._abc_6362_n3558_1), .Y(dp.rf._abc_6362_n3506) );
	NAND2X1 NAND2X1_2038 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3560_1) );
	NAND2X1 NAND2X1_2039 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<29>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3561_1) );
	NAND2X1 NAND2X1_2040 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3560_1), .B(dp.rf._abc_6362_n3561_1), .Y(dp.rf._abc_6362_n3507) );
	NAND2X1 NAND2X1_2041 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3563_1) );
	NAND2X1 NAND2X1_2042 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<30>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3564_1) );
	NAND2X1 NAND2X1_2043 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3563_1), .B(dp.rf._abc_6362_n3564_1), .Y(dp.rf._abc_6362_n3508) );
	NAND2X1 NAND2X1_2044 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n3471_1), .Y(dp.rf._abc_6362_n3566_1) );
	NAND2X1 NAND2X1_2045 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_21_<31>), .B(dp.rf._abc_6362_n3473_1), .Y(dp.rf._abc_6362_n3567_1) );
	NAND2X1 NAND2X1_2046 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3566_1), .B(dp.rf._abc_6362_n3567_1), .Y(dp.rf._abc_6362_n3509) );
	NOR2X1 NOR2X1_205 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2272), .B(dp.rf._abc_6362_n3369_1), .Y(dp.rf._abc_6362_n3569_1) );
	INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3569_1), .Y(dp.rf._abc_6362_n3570_1) );
	NOR2X1 NOR2X1_206 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n3570_1), .Y(dp.rf._abc_6362_n3571_1) );
	NAND2X1 NAND2X1_2047 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3572_1) );
	INVX8 INVX8_19 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3573_1) );
	NAND2X1 NAND2X1_2048 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<0>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3574_1) );
	NAND2X1 NAND2X1_2049 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3572_1), .B(dp.rf._abc_6362_n3574_1), .Y(dp.rf._abc_6362_n3510) );
	NAND2X1 NAND2X1_2050 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3576_1) );
	NAND2X1 NAND2X1_2051 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<1>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3577_1) );
	NAND2X1 NAND2X1_2052 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3576_1), .B(dp.rf._abc_6362_n3577_1), .Y(dp.rf._abc_6362_n3511) );
	NAND2X1 NAND2X1_2053 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3579_1) );
	NAND2X1 NAND2X1_2054 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<2>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3580_1) );
	NAND2X1 NAND2X1_2055 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3579_1), .B(dp.rf._abc_6362_n3580_1), .Y(dp.rf._abc_6362_n3512) );
	NAND2X1 NAND2X1_2056 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3582_1) );
	NAND2X1 NAND2X1_2057 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<3>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3583_1) );
	NAND2X1 NAND2X1_2058 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3582_1), .B(dp.rf._abc_6362_n3583_1), .Y(dp.rf._abc_6362_n3513) );
	NAND2X1 NAND2X1_2059 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3585_1) );
	NAND2X1 NAND2X1_2060 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<4>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3586_1) );
	NAND2X1 NAND2X1_2061 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3585_1), .B(dp.rf._abc_6362_n3586_1), .Y(dp.rf._abc_6362_n3514) );
	NAND2X1 NAND2X1_2062 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3588_1) );
	NAND2X1 NAND2X1_2063 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<5>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3589_1) );
	NAND2X1 NAND2X1_2064 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3588_1), .B(dp.rf._abc_6362_n3589_1), .Y(dp.rf._abc_6362_n3515) );
	NAND2X1 NAND2X1_2065 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3591_1) );
	NAND2X1 NAND2X1_2066 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<6>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3592_1) );
	NAND2X1 NAND2X1_2067 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3591_1), .B(dp.rf._abc_6362_n3592_1), .Y(dp.rf._abc_6362_n3516) );
	NAND2X1 NAND2X1_2068 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3594_1) );
	NAND2X1 NAND2X1_2069 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<7>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3595_1) );
	NAND2X1 NAND2X1_2070 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3594_1), .B(dp.rf._abc_6362_n3595_1), .Y(dp.rf._abc_6362_n3517) );
	NAND2X1 NAND2X1_2071 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3597_1) );
	NAND2X1 NAND2X1_2072 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<8>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3598_1) );
	NAND2X1 NAND2X1_2073 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3597_1), .B(dp.rf._abc_6362_n3598_1), .Y(dp.rf._abc_6362_n3518) );
	NAND2X1 NAND2X1_2074 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3600_1) );
	NAND2X1 NAND2X1_2075 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<9>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3601_1) );
	NAND2X1 NAND2X1_2076 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3600_1), .B(dp.rf._abc_6362_n3601_1), .Y(dp.rf._abc_6362_n3519) );
	NAND2X1 NAND2X1_2077 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3603_1) );
	NAND2X1 NAND2X1_2078 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<10>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3604_1) );
	NAND2X1 NAND2X1_2079 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3603_1), .B(dp.rf._abc_6362_n3604_1), .Y(dp.rf._abc_6362_n3520) );
	NAND2X1 NAND2X1_2080 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3606_1) );
	NAND2X1 NAND2X1_2081 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<11>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3607_1) );
	NAND2X1 NAND2X1_2082 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3606_1), .B(dp.rf._abc_6362_n3607_1), .Y(dp.rf._abc_6362_n3521) );
	NAND2X1 NAND2X1_2083 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3609_1) );
	NAND2X1 NAND2X1_2084 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<12>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3610_1) );
	NAND2X1 NAND2X1_2085 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3609_1), .B(dp.rf._abc_6362_n3610_1), .Y(dp.rf._abc_6362_n3522) );
	NAND2X1 NAND2X1_2086 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3612_1) );
	NAND2X1 NAND2X1_2087 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<13>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3613_1) );
	NAND2X1 NAND2X1_2088 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3612_1), .B(dp.rf._abc_6362_n3613_1), .Y(dp.rf._abc_6362_n3523) );
	NAND2X1 NAND2X1_2089 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3615_1) );
	NAND2X1 NAND2X1_2090 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<14>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3616_1) );
	NAND2X1 NAND2X1_2091 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3615_1), .B(dp.rf._abc_6362_n3616_1), .Y(dp.rf._abc_6362_n3524) );
	NAND2X1 NAND2X1_2092 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3618_1) );
	NAND2X1 NAND2X1_2093 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<15>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3619_1) );
	NAND2X1 NAND2X1_2094 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3618_1), .B(dp.rf._abc_6362_n3619_1), .Y(dp.rf._abc_6362_n3525) );
	NAND2X1 NAND2X1_2095 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3621_1) );
	NAND2X1 NAND2X1_2096 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<16>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3622_1) );
	NAND2X1 NAND2X1_2097 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3621_1), .B(dp.rf._abc_6362_n3622_1), .Y(dp.rf._abc_6362_n3526) );
	NAND2X1 NAND2X1_2098 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3624_1) );
	NAND2X1 NAND2X1_2099 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<17>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3625_1) );
	NAND2X1 NAND2X1_2100 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3624_1), .B(dp.rf._abc_6362_n3625_1), .Y(dp.rf._abc_6362_n3527) );
	NAND2X1 NAND2X1_2101 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3627_1) );
	NAND2X1 NAND2X1_2102 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<18>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3628_1) );
	NAND2X1 NAND2X1_2103 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3627_1), .B(dp.rf._abc_6362_n3628_1), .Y(dp.rf._abc_6362_n3528) );
	NAND2X1 NAND2X1_2104 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3630_1) );
	NAND2X1 NAND2X1_2105 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<19>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3631_1) );
	NAND2X1 NAND2X1_2106 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3630_1), .B(dp.rf._abc_6362_n3631_1), .Y(dp.rf._abc_6362_n3529) );
	NAND2X1 NAND2X1_2107 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3633_1) );
	NAND2X1 NAND2X1_2108 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<20>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3634_1) );
	NAND2X1 NAND2X1_2109 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3633_1), .B(dp.rf._abc_6362_n3634_1), .Y(dp.rf._abc_6362_n3530) );
	NAND2X1 NAND2X1_2110 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3636_1) );
	NAND2X1 NAND2X1_2111 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<21>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3637_1) );
	NAND2X1 NAND2X1_2112 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3636_1), .B(dp.rf._abc_6362_n3637_1), .Y(dp.rf._abc_6362_n3531) );
	NAND2X1 NAND2X1_2113 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3639_1) );
	NAND2X1 NAND2X1_2114 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<22>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3640_1) );
	NAND2X1 NAND2X1_2115 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3639_1), .B(dp.rf._abc_6362_n3640_1), .Y(dp.rf._abc_6362_n3532) );
	NAND2X1 NAND2X1_2116 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3642_1) );
	NAND2X1 NAND2X1_2117 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<23>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3643_1) );
	NAND2X1 NAND2X1_2118 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3642_1), .B(dp.rf._abc_6362_n3643_1), .Y(dp.rf._abc_6362_n3533) );
	NAND2X1 NAND2X1_2119 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3645_1) );
	NAND2X1 NAND2X1_2120 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<24>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3646_1) );
	NAND2X1 NAND2X1_2121 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3645_1), .B(dp.rf._abc_6362_n3646_1), .Y(dp.rf._abc_6362_n3534) );
	NAND2X1 NAND2X1_2122 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3648_1) );
	NAND2X1 NAND2X1_2123 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<25>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3649_1) );
	NAND2X1 NAND2X1_2124 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3648_1), .B(dp.rf._abc_6362_n3649_1), .Y(dp.rf._abc_6362_n3535) );
	NAND2X1 NAND2X1_2125 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3651_1) );
	NAND2X1 NAND2X1_2126 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<26>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3652_1) );
	NAND2X1 NAND2X1_2127 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3651_1), .B(dp.rf._abc_6362_n3652_1), .Y(dp.rf._abc_6362_n3536) );
	NAND2X1 NAND2X1_2128 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3654_1) );
	NAND2X1 NAND2X1_2129 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<27>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3655_1) );
	NAND2X1 NAND2X1_2130 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3654_1), .B(dp.rf._abc_6362_n3655_1), .Y(dp.rf._abc_6362_n3537) );
	NAND2X1 NAND2X1_2131 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3657_1) );
	NAND2X1 NAND2X1_2132 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<28>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3658_1) );
	NAND2X1 NAND2X1_2133 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3657_1), .B(dp.rf._abc_6362_n3658_1), .Y(dp.rf._abc_6362_n3538) );
	NAND2X1 NAND2X1_2134 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3660_1) );
	NAND2X1 NAND2X1_2135 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<29>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3661_1) );
	NAND2X1 NAND2X1_2136 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3660_1), .B(dp.rf._abc_6362_n3661_1), .Y(dp.rf._abc_6362_n3539) );
	NAND2X1 NAND2X1_2137 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3663_1) );
	NAND2X1 NAND2X1_2138 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<30>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3664_1) );
	NAND2X1 NAND2X1_2139 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3663_1), .B(dp.rf._abc_6362_n3664_1), .Y(dp.rf._abc_6362_n3540) );
	NAND2X1 NAND2X1_2140 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n3571_1), .Y(dp.rf._abc_6362_n3666_1) );
	NAND2X1 NAND2X1_2141 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<31>), .B(dp.rf._abc_6362_n3573_1), .Y(dp.rf._abc_6362_n3667_1) );
	NAND2X1 NAND2X1_2142 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3666_1), .B(dp.rf._abc_6362_n3667_1), .Y(dp.rf._abc_6362_n3541) );
	NAND2X1 NAND2X1_2143 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3370_1), .B(dp.rf._abc_6362_n2376), .Y(dp.rf._abc_6362_n3669_1) );
	NOR2X1 NOR2X1_207 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n3669_1), .Y(dp.rf._abc_6362_n3670_1) );
	NAND2X1 NAND2X1_2144 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3671_1) );
	INVX8 INVX8_20 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3672_1) );
	NAND2X1 NAND2X1_2145 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<0>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3673_1) );
	NAND2X1 NAND2X1_2146 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3671_1), .B(dp.rf._abc_6362_n3673_1), .Y(dp.rf._abc_6362_n3542) );
	NAND2X1 NAND2X1_2147 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3675_1) );
	NAND2X1 NAND2X1_2148 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<1>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3676_1) );
	NAND2X1 NAND2X1_2149 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3675_1), .B(dp.rf._abc_6362_n3676_1), .Y(dp.rf._abc_6362_n3543) );
	NAND2X1 NAND2X1_2150 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3678_1) );
	NAND2X1 NAND2X1_2151 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<2>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3679_1) );
	NAND2X1 NAND2X1_2152 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3678_1), .B(dp.rf._abc_6362_n3679_1), .Y(dp.rf._abc_6362_n3544) );
	NAND2X1 NAND2X1_2153 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3681_1) );
	NAND2X1 NAND2X1_2154 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<3>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3682_1) );
	NAND2X1 NAND2X1_2155 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3681_1), .B(dp.rf._abc_6362_n3682_1), .Y(dp.rf._abc_6362_n3545) );
	NAND2X1 NAND2X1_2156 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3684_1) );
	NAND2X1 NAND2X1_2157 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<4>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3685_1) );
	NAND2X1 NAND2X1_2158 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3684_1), .B(dp.rf._abc_6362_n3685_1), .Y(dp.rf._abc_6362_n3546) );
	NAND2X1 NAND2X1_2159 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3687_1) );
	NAND2X1 NAND2X1_2160 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<5>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3688_1) );
	NAND2X1 NAND2X1_2161 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3687_1), .B(dp.rf._abc_6362_n3688_1), .Y(dp.rf._abc_6362_n3547) );
	NAND2X1 NAND2X1_2162 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3690_1) );
	NAND2X1 NAND2X1_2163 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<6>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3691_1) );
	NAND2X1 NAND2X1_2164 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3690_1), .B(dp.rf._abc_6362_n3691_1), .Y(dp.rf._abc_6362_n3548) );
	NAND2X1 NAND2X1_2165 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3693_1) );
	NAND2X1 NAND2X1_2166 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<7>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3694_1) );
	NAND2X1 NAND2X1_2167 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3693_1), .B(dp.rf._abc_6362_n3694_1), .Y(dp.rf._abc_6362_n3549) );
	NAND2X1 NAND2X1_2168 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3696_1) );
	NAND2X1 NAND2X1_2169 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<8>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3697_1) );
	NAND2X1 NAND2X1_2170 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3696_1), .B(dp.rf._abc_6362_n3697_1), .Y(dp.rf._abc_6362_n3550) );
	NAND2X1 NAND2X1_2171 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3699_1) );
	NAND2X1 NAND2X1_2172 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<9>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3700_1) );
	NAND2X1 NAND2X1_2173 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3699_1), .B(dp.rf._abc_6362_n3700_1), .Y(dp.rf._abc_6362_n3551) );
	NAND2X1 NAND2X1_2174 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3702_1) );
	NAND2X1 NAND2X1_2175 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<10>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3703_1) );
	NAND2X1 NAND2X1_2176 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3702_1), .B(dp.rf._abc_6362_n3703_1), .Y(dp.rf._abc_6362_n3552) );
	NAND2X1 NAND2X1_2177 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3705_1) );
	NAND2X1 NAND2X1_2178 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<11>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3706_1) );
	NAND2X1 NAND2X1_2179 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3705_1), .B(dp.rf._abc_6362_n3706_1), .Y(dp.rf._abc_6362_n3553) );
	NAND2X1 NAND2X1_2180 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3708_1) );
	NAND2X1 NAND2X1_2181 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<12>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3709_1) );
	NAND2X1 NAND2X1_2182 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3708_1), .B(dp.rf._abc_6362_n3709_1), .Y(dp.rf._abc_6362_n3554) );
	NAND2X1 NAND2X1_2183 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3711_1) );
	NAND2X1 NAND2X1_2184 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<13>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3712_1) );
	NAND2X1 NAND2X1_2185 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3711_1), .B(dp.rf._abc_6362_n3712_1), .Y(dp.rf._abc_6362_n3555) );
	NAND2X1 NAND2X1_2186 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3714_1) );
	NAND2X1 NAND2X1_2187 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<14>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3715_1) );
	NAND2X1 NAND2X1_2188 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3714_1), .B(dp.rf._abc_6362_n3715_1), .Y(dp.rf._abc_6362_n3556) );
	NAND2X1 NAND2X1_2189 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3717_1) );
	NAND2X1 NAND2X1_2190 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<15>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3718_1) );
	NAND2X1 NAND2X1_2191 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3717_1), .B(dp.rf._abc_6362_n3718_1), .Y(dp.rf._abc_6362_n3557) );
	NAND2X1 NAND2X1_2192 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3720_1) );
	NAND2X1 NAND2X1_2193 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<16>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3721_1) );
	NAND2X1 NAND2X1_2194 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3720_1), .B(dp.rf._abc_6362_n3721_1), .Y(dp.rf._abc_6362_n3558) );
	NAND2X1 NAND2X1_2195 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3723_1) );
	NAND2X1 NAND2X1_2196 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<17>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3724_1) );
	NAND2X1 NAND2X1_2197 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3723_1), .B(dp.rf._abc_6362_n3724_1), .Y(dp.rf._abc_6362_n3559) );
	NAND2X1 NAND2X1_2198 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3726_1) );
	NAND2X1 NAND2X1_2199 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<18>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3727_1) );
	NAND2X1 NAND2X1_2200 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3726_1), .B(dp.rf._abc_6362_n3727_1), .Y(dp.rf._abc_6362_n3560) );
	NAND2X1 NAND2X1_2201 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3729_1) );
	NAND2X1 NAND2X1_2202 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<19>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3730_1) );
	NAND2X1 NAND2X1_2203 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3729_1), .B(dp.rf._abc_6362_n3730_1), .Y(dp.rf._abc_6362_n3561) );
	NAND2X1 NAND2X1_2204 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3732_1) );
	NAND2X1 NAND2X1_2205 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<20>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3733_1) );
	NAND2X1 NAND2X1_2206 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3732_1), .B(dp.rf._abc_6362_n3733_1), .Y(dp.rf._abc_6362_n3562) );
	NAND2X1 NAND2X1_2207 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3735_1) );
	NAND2X1 NAND2X1_2208 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<21>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3736_1) );
	NAND2X1 NAND2X1_2209 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3735_1), .B(dp.rf._abc_6362_n3736_1), .Y(dp.rf._abc_6362_n3563) );
	NAND2X1 NAND2X1_2210 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3738_1) );
	NAND2X1 NAND2X1_2211 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<22>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3739_1) );
	NAND2X1 NAND2X1_2212 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3738_1), .B(dp.rf._abc_6362_n3739_1), .Y(dp.rf._abc_6362_n3564) );
	NAND2X1 NAND2X1_2213 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3741_1) );
	NAND2X1 NAND2X1_2214 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<23>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3742_1) );
	NAND2X1 NAND2X1_2215 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3741_1), .B(dp.rf._abc_6362_n3742_1), .Y(dp.rf._abc_6362_n3565) );
	NAND2X1 NAND2X1_2216 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3744_1) );
	NAND2X1 NAND2X1_2217 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<24>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3745_1) );
	NAND2X1 NAND2X1_2218 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3744_1), .B(dp.rf._abc_6362_n3745_1), .Y(dp.rf._abc_6362_n3566) );
	NAND2X1 NAND2X1_2219 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3747_1) );
	NAND2X1 NAND2X1_2220 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<25>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3748_1) );
	NAND2X1 NAND2X1_2221 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3747_1), .B(dp.rf._abc_6362_n3748_1), .Y(dp.rf._abc_6362_n3567) );
	NAND2X1 NAND2X1_2222 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3750_1) );
	NAND2X1 NAND2X1_2223 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<26>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3751_1) );
	NAND2X1 NAND2X1_2224 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3750_1), .B(dp.rf._abc_6362_n3751_1), .Y(dp.rf._abc_6362_n3568) );
	NAND2X1 NAND2X1_2225 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3753_1) );
	NAND2X1 NAND2X1_2226 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<27>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3754_1) );
	NAND2X1 NAND2X1_2227 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3753_1), .B(dp.rf._abc_6362_n3754_1), .Y(dp.rf._abc_6362_n3569) );
	NAND2X1 NAND2X1_2228 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3756_1) );
	NAND2X1 NAND2X1_2229 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<28>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3757_1) );
	NAND2X1 NAND2X1_2230 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3756_1), .B(dp.rf._abc_6362_n3757_1), .Y(dp.rf._abc_6362_n3570) );
	NAND2X1 NAND2X1_2231 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3759_1) );
	NAND2X1 NAND2X1_2232 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<29>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3760_1) );
	NAND2X1 NAND2X1_2233 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3759_1), .B(dp.rf._abc_6362_n3760_1), .Y(dp.rf._abc_6362_n3571) );
	NAND2X1 NAND2X1_2234 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3762_1) );
	NAND2X1 NAND2X1_2235 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<30>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3763_1) );
	NAND2X1 NAND2X1_2236 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3762_1), .B(dp.rf._abc_6362_n3763_1), .Y(dp.rf._abc_6362_n3572) );
	NAND2X1 NAND2X1_2237 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n3670_1), .Y(dp.rf._abc_6362_n3765_1) );
	NAND2X1 NAND2X1_2238 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_23_<31>), .B(dp.rf._abc_6362_n3672_1), .Y(dp.rf._abc_6362_n3766_1) );
	NAND2X1 NAND2X1_2239 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3765_1), .B(dp.rf._abc_6362_n3766_1), .Y(dp.rf._abc_6362_n3573) );
	NAND2X1 NAND2X1_2240 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2167), .B(dp.rf._abc_6362_n2275), .Y(dp.rf._abc_6362_n3768_1) );
	NOR2X1 NOR2X1_208 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n3768_1), .Y(dp.rf._abc_6362_n3769_1) );
	NAND2X1 NAND2X1_2241 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3770_1) );
	INVX8 INVX8_21 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3771_1) );
	NAND2X1 NAND2X1_2242 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<0>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3772_1) );
	NAND2X1 NAND2X1_2243 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3770_1), .B(dp.rf._abc_6362_n3772_1), .Y(dp.rf._abc_6362_n3574) );
	NAND2X1 NAND2X1_2244 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3774_1) );
	NAND2X1 NAND2X1_2245 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<1>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3775_1) );
	NAND2X1 NAND2X1_2246 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3774_1), .B(dp.rf._abc_6362_n3775_1), .Y(dp.rf._abc_6362_n3575) );
	NAND2X1 NAND2X1_2247 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3777_1) );
	NAND2X1 NAND2X1_2248 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<2>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3778_1) );
	NAND2X1 NAND2X1_2249 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3777_1), .B(dp.rf._abc_6362_n3778_1), .Y(dp.rf._abc_6362_n3576) );
	NAND2X1 NAND2X1_2250 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3780_1) );
	NAND2X1 NAND2X1_2251 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<3>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3781_1) );
	NAND2X1 NAND2X1_2252 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3780_1), .B(dp.rf._abc_6362_n3781_1), .Y(dp.rf._abc_6362_n3577) );
	NAND2X1 NAND2X1_2253 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3783_1) );
	NAND2X1 NAND2X1_2254 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<4>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3784_1) );
	NAND2X1 NAND2X1_2255 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3783_1), .B(dp.rf._abc_6362_n3784_1), .Y(dp.rf._abc_6362_n3578) );
	NAND2X1 NAND2X1_2256 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3786_1) );
	NAND2X1 NAND2X1_2257 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<5>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3787_1) );
	NAND2X1 NAND2X1_2258 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3786_1), .B(dp.rf._abc_6362_n3787_1), .Y(dp.rf._abc_6362_n3579) );
	NAND2X1 NAND2X1_2259 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3789_1) );
	NAND2X1 NAND2X1_2260 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<6>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3790_1) );
	NAND2X1 NAND2X1_2261 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3789_1), .B(dp.rf._abc_6362_n3790_1), .Y(dp.rf._abc_6362_n3580) );
	NAND2X1 NAND2X1_2262 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3792_1) );
	NAND2X1 NAND2X1_2263 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<7>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3793_1) );
	NAND2X1 NAND2X1_2264 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3792_1), .B(dp.rf._abc_6362_n3793_1), .Y(dp.rf._abc_6362_n3581) );
	NAND2X1 NAND2X1_2265 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3795_1) );
	NAND2X1 NAND2X1_2266 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<8>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3796_1) );
	NAND2X1 NAND2X1_2267 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3795_1), .B(dp.rf._abc_6362_n3796_1), .Y(dp.rf._abc_6362_n3582) );
	NAND2X1 NAND2X1_2268 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3798_1) );
	NAND2X1 NAND2X1_2269 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<9>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3799_1) );
	NAND2X1 NAND2X1_2270 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3798_1), .B(dp.rf._abc_6362_n3799_1), .Y(dp.rf._abc_6362_n3583) );
	NAND2X1 NAND2X1_2271 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3801_1) );
	NAND2X1 NAND2X1_2272 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<10>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3802_1) );
	NAND2X1 NAND2X1_2273 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3801_1), .B(dp.rf._abc_6362_n3802_1), .Y(dp.rf._abc_6362_n3584) );
	NAND2X1 NAND2X1_2274 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3804_1) );
	NAND2X1 NAND2X1_2275 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<11>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3805_1) );
	NAND2X1 NAND2X1_2276 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3804_1), .B(dp.rf._abc_6362_n3805_1), .Y(dp.rf._abc_6362_n3585) );
	NAND2X1 NAND2X1_2277 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3807_1) );
	NAND2X1 NAND2X1_2278 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<12>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3808_1) );
	NAND2X1 NAND2X1_2279 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3807_1), .B(dp.rf._abc_6362_n3808_1), .Y(dp.rf._abc_6362_n3586) );
	NAND2X1 NAND2X1_2280 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3810_1) );
	NAND2X1 NAND2X1_2281 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<13>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3811_1) );
	NAND2X1 NAND2X1_2282 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3810_1), .B(dp.rf._abc_6362_n3811_1), .Y(dp.rf._abc_6362_n3587) );
	NAND2X1 NAND2X1_2283 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3813_1) );
	NAND2X1 NAND2X1_2284 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<14>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3814_1) );
	NAND2X1 NAND2X1_2285 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3813_1), .B(dp.rf._abc_6362_n3814_1), .Y(dp.rf._abc_6362_n3588) );
	NAND2X1 NAND2X1_2286 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3816_1) );
	NAND2X1 NAND2X1_2287 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<15>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3817_1) );
	NAND2X1 NAND2X1_2288 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3816_1), .B(dp.rf._abc_6362_n3817_1), .Y(dp.rf._abc_6362_n3589) );
	NAND2X1 NAND2X1_2289 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3819_1) );
	NAND2X1 NAND2X1_2290 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<16>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3820_1) );
	NAND2X1 NAND2X1_2291 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3819_1), .B(dp.rf._abc_6362_n3820_1), .Y(dp.rf._abc_6362_n3590) );
	NAND2X1 NAND2X1_2292 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3822_1) );
	NAND2X1 NAND2X1_2293 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<17>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3823_1) );
	NAND2X1 NAND2X1_2294 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3822_1), .B(dp.rf._abc_6362_n3823_1), .Y(dp.rf._abc_6362_n3591) );
	NAND2X1 NAND2X1_2295 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3825_1) );
	NAND2X1 NAND2X1_2296 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<18>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3826_1) );
	NAND2X1 NAND2X1_2297 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3825_1), .B(dp.rf._abc_6362_n3826_1), .Y(dp.rf._abc_6362_n3592) );
	NAND2X1 NAND2X1_2298 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3828_1) );
	NAND2X1 NAND2X1_2299 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<19>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3829_1) );
	NAND2X1 NAND2X1_2300 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3828_1), .B(dp.rf._abc_6362_n3829_1), .Y(dp.rf._abc_6362_n3593) );
	NAND2X1 NAND2X1_2301 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3831_1) );
	NAND2X1 NAND2X1_2302 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<20>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3832_1) );
	NAND2X1 NAND2X1_2303 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3831_1), .B(dp.rf._abc_6362_n3832_1), .Y(dp.rf._abc_6362_n3594) );
	NAND2X1 NAND2X1_2304 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3834_1) );
	NAND2X1 NAND2X1_2305 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<21>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3835_1) );
	NAND2X1 NAND2X1_2306 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3834_1), .B(dp.rf._abc_6362_n3835_1), .Y(dp.rf._abc_6362_n3595) );
	NAND2X1 NAND2X1_2307 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3837_1) );
	NAND2X1 NAND2X1_2308 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<22>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3838_1) );
	NAND2X1 NAND2X1_2309 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3837_1), .B(dp.rf._abc_6362_n3838_1), .Y(dp.rf._abc_6362_n3596) );
	NAND2X1 NAND2X1_2310 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3840_1) );
	NAND2X1 NAND2X1_2311 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<23>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3841_1) );
	NAND2X1 NAND2X1_2312 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3840_1), .B(dp.rf._abc_6362_n3841_1), .Y(dp.rf._abc_6362_n3597) );
	NAND2X1 NAND2X1_2313 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3843_1) );
	NAND2X1 NAND2X1_2314 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<24>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3844_1) );
	NAND2X1 NAND2X1_2315 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3843_1), .B(dp.rf._abc_6362_n3844_1), .Y(dp.rf._abc_6362_n3598) );
	NAND2X1 NAND2X1_2316 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3846_1) );
	NAND2X1 NAND2X1_2317 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<25>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3847_1) );
	NAND2X1 NAND2X1_2318 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3846_1), .B(dp.rf._abc_6362_n3847_1), .Y(dp.rf._abc_6362_n3599) );
	NAND2X1 NAND2X1_2319 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3849_1) );
	NAND2X1 NAND2X1_2320 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<26>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3850_1) );
	NAND2X1 NAND2X1_2321 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3849_1), .B(dp.rf._abc_6362_n3850_1), .Y(dp.rf._abc_6362_n3600) );
	NAND2X1 NAND2X1_2322 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3852_1) );
	NAND2X1 NAND2X1_2323 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<27>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3853_1) );
	NAND2X1 NAND2X1_2324 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3852_1), .B(dp.rf._abc_6362_n3853_1), .Y(dp.rf._abc_6362_n3601) );
	NAND2X1 NAND2X1_2325 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3855_1) );
	NAND2X1 NAND2X1_2326 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<28>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3856_1) );
	NAND2X1 NAND2X1_2327 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3855_1), .B(dp.rf._abc_6362_n3856_1), .Y(dp.rf._abc_6362_n3602) );
	NAND2X1 NAND2X1_2328 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3858_1) );
	NAND2X1 NAND2X1_2329 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<29>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3859_1) );
	NAND2X1 NAND2X1_2330 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3858_1), .B(dp.rf._abc_6362_n3859_1), .Y(dp.rf._abc_6362_n3603) );
	NAND2X1 NAND2X1_2331 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3861_1) );
	NAND2X1 NAND2X1_2332 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<30>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3862_1) );
	NAND2X1 NAND2X1_2333 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3861_1), .B(dp.rf._abc_6362_n3862_1), .Y(dp.rf._abc_6362_n3604) );
	NAND2X1 NAND2X1_2334 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n3769_1), .Y(dp.rf._abc_6362_n3864_1) );
	NAND2X1 NAND2X1_2335 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<31>), .B(dp.rf._abc_6362_n3771_1), .Y(dp.rf._abc_6362_n3865_1) );
	NAND2X1 NAND2X1_2336 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3864_1), .B(dp.rf._abc_6362_n3865_1), .Y(dp.rf._abc_6362_n3605) );
	NAND2X1 NAND2X1_2337 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2275), .B(dp.rf._abc_6362_n2576), .Y(dp.rf._abc_6362_n3867_1) );
	NOR2X1 NOR2X1_209 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n3867_1), .Y(dp.rf._abc_6362_n3868_1) );
	NAND2X1 NAND2X1_2338 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3869_1) );
	INVX8 INVX8_22 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3870_1) );
	NAND2X1 NAND2X1_2339 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<0>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3871_1) );
	NAND2X1 NAND2X1_2340 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3869_1), .B(dp.rf._abc_6362_n3871_1), .Y(dp.rf._abc_6362_n3606) );
	NAND2X1 NAND2X1_2341 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3873_1) );
	NAND2X1 NAND2X1_2342 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<1>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3874_1) );
	NAND2X1 NAND2X1_2343 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3873_1), .B(dp.rf._abc_6362_n3874_1), .Y(dp.rf._abc_6362_n3607) );
	NAND2X1 NAND2X1_2344 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3876_1) );
	NAND2X1 NAND2X1_2345 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<2>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3877_1) );
	NAND2X1 NAND2X1_2346 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3876_1), .B(dp.rf._abc_6362_n3877_1), .Y(dp.rf._abc_6362_n3608) );
	NAND2X1 NAND2X1_2347 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3879_1) );
	NAND2X1 NAND2X1_2348 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<3>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3880_1) );
	NAND2X1 NAND2X1_2349 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3879_1), .B(dp.rf._abc_6362_n3880_1), .Y(dp.rf._abc_6362_n3609) );
	NAND2X1 NAND2X1_2350 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3882_1) );
	NAND2X1 NAND2X1_2351 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<4>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3883_1) );
	NAND2X1 NAND2X1_2352 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3882_1), .B(dp.rf._abc_6362_n3883_1), .Y(dp.rf._abc_6362_n3610) );
	NAND2X1 NAND2X1_2353 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3885_1) );
	NAND2X1 NAND2X1_2354 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<5>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3886_1) );
	NAND2X1 NAND2X1_2355 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3885_1), .B(dp.rf._abc_6362_n3886_1), .Y(dp.rf._abc_6362_n3611) );
	NAND2X1 NAND2X1_2356 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3888_1) );
	NAND2X1 NAND2X1_2357 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<6>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3889_1) );
	NAND2X1 NAND2X1_2358 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3888_1), .B(dp.rf._abc_6362_n3889_1), .Y(dp.rf._abc_6362_n3612) );
	NAND2X1 NAND2X1_2359 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3891_1) );
	NAND2X1 NAND2X1_2360 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<7>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3892_1) );
	NAND2X1 NAND2X1_2361 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3891_1), .B(dp.rf._abc_6362_n3892_1), .Y(dp.rf._abc_6362_n3613) );
	NAND2X1 NAND2X1_2362 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3894_1) );
	NAND2X1 NAND2X1_2363 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<8>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3895_1) );
	NAND2X1 NAND2X1_2364 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3894_1), .B(dp.rf._abc_6362_n3895_1), .Y(dp.rf._abc_6362_n3614) );
	NAND2X1 NAND2X1_2365 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3897_1) );
	NAND2X1 NAND2X1_2366 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<9>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3898_1) );
	NAND2X1 NAND2X1_2367 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3897_1), .B(dp.rf._abc_6362_n3898_1), .Y(dp.rf._abc_6362_n3615) );
	NAND2X1 NAND2X1_2368 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3900_1) );
	NAND2X1 NAND2X1_2369 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<10>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3901_1) );
	NAND2X1 NAND2X1_2370 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3900_1), .B(dp.rf._abc_6362_n3901_1), .Y(dp.rf._abc_6362_n3616) );
	NAND2X1 NAND2X1_2371 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3903_1) );
	NAND2X1 NAND2X1_2372 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<11>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3904_1) );
	NAND2X1 NAND2X1_2373 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3903_1), .B(dp.rf._abc_6362_n3904_1), .Y(dp.rf._abc_6362_n3617) );
	NAND2X1 NAND2X1_2374 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3906_1) );
	NAND2X1 NAND2X1_2375 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<12>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3907_1) );
	NAND2X1 NAND2X1_2376 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3906_1), .B(dp.rf._abc_6362_n3907_1), .Y(dp.rf._abc_6362_n3618) );
	NAND2X1 NAND2X1_2377 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3909_1) );
	NAND2X1 NAND2X1_2378 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<13>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3910_1) );
	NAND2X1 NAND2X1_2379 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3909_1), .B(dp.rf._abc_6362_n3910_1), .Y(dp.rf._abc_6362_n3619) );
	NAND2X1 NAND2X1_2380 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3912_1) );
	NAND2X1 NAND2X1_2381 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<14>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3913_1) );
	NAND2X1 NAND2X1_2382 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3912_1), .B(dp.rf._abc_6362_n3913_1), .Y(dp.rf._abc_6362_n3620) );
	NAND2X1 NAND2X1_2383 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3915_1) );
	NAND2X1 NAND2X1_2384 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<15>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3916_1) );
	NAND2X1 NAND2X1_2385 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3915_1), .B(dp.rf._abc_6362_n3916_1), .Y(dp.rf._abc_6362_n3621) );
	NAND2X1 NAND2X1_2386 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3918_1) );
	NAND2X1 NAND2X1_2387 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<16>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3919_1) );
	NAND2X1 NAND2X1_2388 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3918_1), .B(dp.rf._abc_6362_n3919_1), .Y(dp.rf._abc_6362_n3622) );
	NAND2X1 NAND2X1_2389 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3921_1) );
	NAND2X1 NAND2X1_2390 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<17>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3922_1) );
	NAND2X1 NAND2X1_2391 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3921_1), .B(dp.rf._abc_6362_n3922_1), .Y(dp.rf._abc_6362_n3623) );
	NAND2X1 NAND2X1_2392 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3924_1) );
	NAND2X1 NAND2X1_2393 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<18>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3925_1) );
	NAND2X1 NAND2X1_2394 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3924_1), .B(dp.rf._abc_6362_n3925_1), .Y(dp.rf._abc_6362_n3624) );
	NAND2X1 NAND2X1_2395 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3927_1) );
	NAND2X1 NAND2X1_2396 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<19>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3928_1) );
	NAND2X1 NAND2X1_2397 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3927_1), .B(dp.rf._abc_6362_n3928_1), .Y(dp.rf._abc_6362_n3625) );
	NAND2X1 NAND2X1_2398 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3930_1) );
	NAND2X1 NAND2X1_2399 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<20>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3931_1) );
	NAND2X1 NAND2X1_2400 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3930_1), .B(dp.rf._abc_6362_n3931_1), .Y(dp.rf._abc_6362_n3626) );
	NAND2X1 NAND2X1_2401 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3933_1) );
	NAND2X1 NAND2X1_2402 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<21>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3934_1) );
	NAND2X1 NAND2X1_2403 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3933_1), .B(dp.rf._abc_6362_n3934_1), .Y(dp.rf._abc_6362_n3627) );
	NAND2X1 NAND2X1_2404 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3936_1) );
	NAND2X1 NAND2X1_2405 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<22>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3937_1) );
	NAND2X1 NAND2X1_2406 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3936_1), .B(dp.rf._abc_6362_n3937_1), .Y(dp.rf._abc_6362_n3628) );
	NAND2X1 NAND2X1_2407 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3939_1) );
	NAND2X1 NAND2X1_2408 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<23>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3940_1) );
	NAND2X1 NAND2X1_2409 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3939_1), .B(dp.rf._abc_6362_n3940_1), .Y(dp.rf._abc_6362_n3629) );
	NAND2X1 NAND2X1_2410 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3942_1) );
	NAND2X1 NAND2X1_2411 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<24>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3943_1) );
	NAND2X1 NAND2X1_2412 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3942_1), .B(dp.rf._abc_6362_n3943_1), .Y(dp.rf._abc_6362_n3630) );
	NAND2X1 NAND2X1_2413 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3945_1) );
	NAND2X1 NAND2X1_2414 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<25>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3946_1) );
	NAND2X1 NAND2X1_2415 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3945_1), .B(dp.rf._abc_6362_n3946_1), .Y(dp.rf._abc_6362_n3631) );
	NAND2X1 NAND2X1_2416 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3948_1) );
	NAND2X1 NAND2X1_2417 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<26>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3949_1) );
	NAND2X1 NAND2X1_2418 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3948_1), .B(dp.rf._abc_6362_n3949_1), .Y(dp.rf._abc_6362_n3632) );
	NAND2X1 NAND2X1_2419 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3951_1) );
	NAND2X1 NAND2X1_2420 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<27>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3952_1) );
	NAND2X1 NAND2X1_2421 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3951_1), .B(dp.rf._abc_6362_n3952_1), .Y(dp.rf._abc_6362_n3633) );
	NAND2X1 NAND2X1_2422 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3954_1) );
	NAND2X1 NAND2X1_2423 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<28>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3955_1) );
	NAND2X1 NAND2X1_2424 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3954_1), .B(dp.rf._abc_6362_n3955_1), .Y(dp.rf._abc_6362_n3634) );
	NAND2X1 NAND2X1_2425 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3957_1) );
	NAND2X1 NAND2X1_2426 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<29>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3958_1) );
	NAND2X1 NAND2X1_2427 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3957_1), .B(dp.rf._abc_6362_n3958_1), .Y(dp.rf._abc_6362_n3635) );
	NAND2X1 NAND2X1_2428 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3960_1) );
	NAND2X1 NAND2X1_2429 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<30>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3961_1) );
	NAND2X1 NAND2X1_2430 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3960_1), .B(dp.rf._abc_6362_n3961_1), .Y(dp.rf._abc_6362_n3636) );
	NAND2X1 NAND2X1_2431 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n3868_1), .Y(dp.rf._abc_6362_n3963_1) );
	NAND2X1 NAND2X1_2432 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_25_<31>), .B(dp.rf._abc_6362_n3870_1), .Y(dp.rf._abc_6362_n3964_1) );
	NAND2X1 NAND2X1_2433 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3963_1), .B(dp.rf._abc_6362_n3964_1), .Y(dp.rf._abc_6362_n3637) );
	NOR2X1 NOR2X1_210 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n2276), .Y(dp.rf._abc_6362_n3966_1) );
	NAND2X1 NAND2X1_2434 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3967_1) );
	INVX8 INVX8_23 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3968_1) );
	NAND2X1 NAND2X1_2435 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<0>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n3969_1) );
	NAND2X1 NAND2X1_2436 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3967_1), .B(dp.rf._abc_6362_n3969_1), .Y(dp.rf._abc_6362_n3638) );
	NAND2X1 NAND2X1_2437 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3971_1) );
	NAND2X1 NAND2X1_2438 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<1>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n3972_1) );
	NAND2X1 NAND2X1_2439 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3971_1), .B(dp.rf._abc_6362_n3972_1), .Y(dp.rf._abc_6362_n3639) );
	NAND2X1 NAND2X1_2440 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3974_1) );
	NAND2X1 NAND2X1_2441 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<2>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n3975_1) );
	NAND2X1 NAND2X1_2442 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3974_1), .B(dp.rf._abc_6362_n3975_1), .Y(dp.rf._abc_6362_n3640) );
	NAND2X1 NAND2X1_2443 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3977_1) );
	NAND2X1 NAND2X1_2444 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<3>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n3978_1) );
	NAND2X1 NAND2X1_2445 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3977_1), .B(dp.rf._abc_6362_n3978_1), .Y(dp.rf._abc_6362_n3641) );
	NAND2X1 NAND2X1_2446 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3980_1) );
	NAND2X1 NAND2X1_2447 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<4>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n3981_1) );
	NAND2X1 NAND2X1_2448 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3980_1), .B(dp.rf._abc_6362_n3981_1), .Y(dp.rf._abc_6362_n3642) );
	NAND2X1 NAND2X1_2449 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3983_1) );
	NAND2X1 NAND2X1_2450 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<5>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n3984_1) );
	NAND2X1 NAND2X1_2451 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3983_1), .B(dp.rf._abc_6362_n3984_1), .Y(dp.rf._abc_6362_n3643) );
	NAND2X1 NAND2X1_2452 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3986_1) );
	NAND2X1 NAND2X1_2453 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<6>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n3987_1) );
	NAND2X1 NAND2X1_2454 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3986_1), .B(dp.rf._abc_6362_n3987_1), .Y(dp.rf._abc_6362_n3644) );
	NAND2X1 NAND2X1_2455 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3989_1) );
	NAND2X1 NAND2X1_2456 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<7>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n3990_1) );
	NAND2X1 NAND2X1_2457 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3989_1), .B(dp.rf._abc_6362_n3990_1), .Y(dp.rf._abc_6362_n3645) );
	NAND2X1 NAND2X1_2458 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3992_1) );
	NAND2X1 NAND2X1_2459 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<8>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n3993_1) );
	NAND2X1 NAND2X1_2460 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3992_1), .B(dp.rf._abc_6362_n3993_1), .Y(dp.rf._abc_6362_n3646) );
	NAND2X1 NAND2X1_2461 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3995_1) );
	NAND2X1 NAND2X1_2462 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<9>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n3996_1) );
	NAND2X1 NAND2X1_2463 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3995_1), .B(dp.rf._abc_6362_n3996_1), .Y(dp.rf._abc_6362_n3647) );
	NAND2X1 NAND2X1_2464 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n3998_1) );
	NAND2X1 NAND2X1_2465 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<10>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n3999_1) );
	NAND2X1 NAND2X1_2466 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n3998_1), .B(dp.rf._abc_6362_n3999_1), .Y(dp.rf._abc_6362_n3648) );
	NAND2X1 NAND2X1_2467 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4001_1) );
	NAND2X1 NAND2X1_2468 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<11>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4002_1) );
	NAND2X1 NAND2X1_2469 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4001_1), .B(dp.rf._abc_6362_n4002_1), .Y(dp.rf._abc_6362_n3649) );
	NAND2X1 NAND2X1_2470 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4004_1) );
	NAND2X1 NAND2X1_2471 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<12>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4005_1) );
	NAND2X1 NAND2X1_2472 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4004_1), .B(dp.rf._abc_6362_n4005_1), .Y(dp.rf._abc_6362_n3650) );
	NAND2X1 NAND2X1_2473 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4007_1) );
	NAND2X1 NAND2X1_2474 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<13>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4008_1) );
	NAND2X1 NAND2X1_2475 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4007_1), .B(dp.rf._abc_6362_n4008_1), .Y(dp.rf._abc_6362_n3651) );
	NAND2X1 NAND2X1_2476 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4010_1) );
	NAND2X1 NAND2X1_2477 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<14>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4011_1) );
	NAND2X1 NAND2X1_2478 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4010_1), .B(dp.rf._abc_6362_n4011_1), .Y(dp.rf._abc_6362_n3652) );
	NAND2X1 NAND2X1_2479 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4013_1) );
	NAND2X1 NAND2X1_2480 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<15>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4014_1) );
	NAND2X1 NAND2X1_2481 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4013_1), .B(dp.rf._abc_6362_n4014_1), .Y(dp.rf._abc_6362_n3653) );
	NAND2X1 NAND2X1_2482 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4016_1) );
	NAND2X1 NAND2X1_2483 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<16>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4017_1) );
	NAND2X1 NAND2X1_2484 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4016_1), .B(dp.rf._abc_6362_n4017_1), .Y(dp.rf._abc_6362_n3654) );
	NAND2X1 NAND2X1_2485 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4019_1) );
	NAND2X1 NAND2X1_2486 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<17>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4020_1) );
	NAND2X1 NAND2X1_2487 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4019_1), .B(dp.rf._abc_6362_n4020_1), .Y(dp.rf._abc_6362_n3655) );
	NAND2X1 NAND2X1_2488 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4022_1) );
	NAND2X1 NAND2X1_2489 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<18>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4023_1) );
	NAND2X1 NAND2X1_2490 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4022_1), .B(dp.rf._abc_6362_n4023_1), .Y(dp.rf._abc_6362_n3656) );
	NAND2X1 NAND2X1_2491 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4025_1) );
	NAND2X1 NAND2X1_2492 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<19>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4026_1) );
	NAND2X1 NAND2X1_2493 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4025_1), .B(dp.rf._abc_6362_n4026_1), .Y(dp.rf._abc_6362_n3657) );
	NAND2X1 NAND2X1_2494 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4028_1) );
	NAND2X1 NAND2X1_2495 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<20>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4029_1) );
	NAND2X1 NAND2X1_2496 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4028_1), .B(dp.rf._abc_6362_n4029_1), .Y(dp.rf._abc_6362_n3658) );
	NAND2X1 NAND2X1_2497 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4031_1) );
	NAND2X1 NAND2X1_2498 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<21>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4032_1) );
	NAND2X1 NAND2X1_2499 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4031_1), .B(dp.rf._abc_6362_n4032_1), .Y(dp.rf._abc_6362_n3659) );
	NAND2X1 NAND2X1_2500 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4034_1) );
	NAND2X1 NAND2X1_2501 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<22>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4035_1) );
	NAND2X1 NAND2X1_2502 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4034_1), .B(dp.rf._abc_6362_n4035_1), .Y(dp.rf._abc_6362_n3660) );
	NAND2X1 NAND2X1_2503 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4037_1) );
	NAND2X1 NAND2X1_2504 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<23>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4038_1) );
	NAND2X1 NAND2X1_2505 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4037_1), .B(dp.rf._abc_6362_n4038_1), .Y(dp.rf._abc_6362_n3661) );
	NAND2X1 NAND2X1_2506 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4040_1) );
	NAND2X1 NAND2X1_2507 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<24>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4041_1) );
	NAND2X1 NAND2X1_2508 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4040_1), .B(dp.rf._abc_6362_n4041_1), .Y(dp.rf._abc_6362_n3662) );
	NAND2X1 NAND2X1_2509 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4043_1) );
	NAND2X1 NAND2X1_2510 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<25>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4044_1) );
	NAND2X1 NAND2X1_2511 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4043_1), .B(dp.rf._abc_6362_n4044_1), .Y(dp.rf._abc_6362_n3663) );
	NAND2X1 NAND2X1_2512 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4046_1) );
	NAND2X1 NAND2X1_2513 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<26>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4047_1) );
	NAND2X1 NAND2X1_2514 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4046_1), .B(dp.rf._abc_6362_n4047_1), .Y(dp.rf._abc_6362_n3664) );
	NAND2X1 NAND2X1_2515 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4049_1) );
	NAND2X1 NAND2X1_2516 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<27>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4050_1) );
	NAND2X1 NAND2X1_2517 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4049_1), .B(dp.rf._abc_6362_n4050_1), .Y(dp.rf._abc_6362_n3665) );
	NAND2X1 NAND2X1_2518 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4052_1) );
	NAND2X1 NAND2X1_2519 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<28>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4053_1) );
	NAND2X1 NAND2X1_2520 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4052_1), .B(dp.rf._abc_6362_n4053_1), .Y(dp.rf._abc_6362_n3666) );
	NAND2X1 NAND2X1_2521 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4055_1) );
	NAND2X1 NAND2X1_2522 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<29>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4056_1) );
	NAND2X1 NAND2X1_2523 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4055_1), .B(dp.rf._abc_6362_n4056_1), .Y(dp.rf._abc_6362_n3667) );
	NAND2X1 NAND2X1_2524 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4058_1) );
	NAND2X1 NAND2X1_2525 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<30>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4059_1) );
	NAND2X1 NAND2X1_2526 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4058_1), .B(dp.rf._abc_6362_n4059_1), .Y(dp.rf._abc_6362_n3668) );
	NAND2X1 NAND2X1_2527 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n3966_1), .Y(dp.rf._abc_6362_n4061_1) );
	NAND2X1 NAND2X1_2528 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<31>), .B(dp.rf._abc_6362_n3968_1), .Y(dp.rf._abc_6362_n4062_1) );
	NAND2X1 NAND2X1_2529 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4061_1), .B(dp.rf._abc_6362_n4062_1), .Y(dp.rf._abc_6362_n3669) );
	NOR2X1 NOR2X1_211 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n2377), .Y(dp.rf._abc_6362_n4064_1) );
	NAND2X1 NAND2X1_2530 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4065_1) );
	INVX8 INVX8_24 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4066_1) );
	NAND2X1 NAND2X1_2531 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<0>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4067_1) );
	NAND2X1 NAND2X1_2532 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4065_1), .B(dp.rf._abc_6362_n4067_1), .Y(dp.rf._abc_6362_n3670) );
	NAND2X1 NAND2X1_2533 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4069_1) );
	NAND2X1 NAND2X1_2534 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<1>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4070_1) );
	NAND2X1 NAND2X1_2535 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4069_1), .B(dp.rf._abc_6362_n4070_1), .Y(dp.rf._abc_6362_n3671) );
	NAND2X1 NAND2X1_2536 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4072_1) );
	NAND2X1 NAND2X1_2537 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<2>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4073_1) );
	NAND2X1 NAND2X1_2538 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4072_1), .B(dp.rf._abc_6362_n4073_1), .Y(dp.rf._abc_6362_n3672) );
	NAND2X1 NAND2X1_2539 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4075_1) );
	NAND2X1 NAND2X1_2540 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<3>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4076_1) );
	NAND2X1 NAND2X1_2541 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4075_1), .B(dp.rf._abc_6362_n4076_1), .Y(dp.rf._abc_6362_n3673) );
	NAND2X1 NAND2X1_2542 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4078_1) );
	NAND2X1 NAND2X1_2543 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<4>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4079_1) );
	NAND2X1 NAND2X1_2544 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4078_1), .B(dp.rf._abc_6362_n4079_1), .Y(dp.rf._abc_6362_n3674) );
	NAND2X1 NAND2X1_2545 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4081_1) );
	NAND2X1 NAND2X1_2546 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<5>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4082_1) );
	NAND2X1 NAND2X1_2547 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4081_1), .B(dp.rf._abc_6362_n4082_1), .Y(dp.rf._abc_6362_n3675) );
	NAND2X1 NAND2X1_2548 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4084_1) );
	NAND2X1 NAND2X1_2549 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<6>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4085_1) );
	NAND2X1 NAND2X1_2550 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4084_1), .B(dp.rf._abc_6362_n4085_1), .Y(dp.rf._abc_6362_n3676) );
	NAND2X1 NAND2X1_2551 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4087_1) );
	NAND2X1 NAND2X1_2552 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<7>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4088_1) );
	NAND2X1 NAND2X1_2553 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4087_1), .B(dp.rf._abc_6362_n4088_1), .Y(dp.rf._abc_6362_n3677) );
	NAND2X1 NAND2X1_2554 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4090_1) );
	NAND2X1 NAND2X1_2555 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<8>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4091_1) );
	NAND2X1 NAND2X1_2556 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4090_1), .B(dp.rf._abc_6362_n4091_1), .Y(dp.rf._abc_6362_n3678) );
	NAND2X1 NAND2X1_2557 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4093_1) );
	NAND2X1 NAND2X1_2558 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<9>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4094_1) );
	NAND2X1 NAND2X1_2559 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4093_1), .B(dp.rf._abc_6362_n4094_1), .Y(dp.rf._abc_6362_n3679) );
	NAND2X1 NAND2X1_2560 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4096_1) );
	NAND2X1 NAND2X1_2561 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<10>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4097_1) );
	NAND2X1 NAND2X1_2562 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4096_1), .B(dp.rf._abc_6362_n4097_1), .Y(dp.rf._abc_6362_n3680) );
	NAND2X1 NAND2X1_2563 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4099_1) );
	NAND2X1 NAND2X1_2564 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<11>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4100_1) );
	NAND2X1 NAND2X1_2565 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4099_1), .B(dp.rf._abc_6362_n4100_1), .Y(dp.rf._abc_6362_n3681) );
	NAND2X1 NAND2X1_2566 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4102_1) );
	NAND2X1 NAND2X1_2567 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<12>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4103_1) );
	NAND2X1 NAND2X1_2568 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4102_1), .B(dp.rf._abc_6362_n4103_1), .Y(dp.rf._abc_6362_n3682) );
	NAND2X1 NAND2X1_2569 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4105_1) );
	NAND2X1 NAND2X1_2570 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<13>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4106_1) );
	NAND2X1 NAND2X1_2571 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4105_1), .B(dp.rf._abc_6362_n4106_1), .Y(dp.rf._abc_6362_n3683) );
	NAND2X1 NAND2X1_2572 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4108_1) );
	NAND2X1 NAND2X1_2573 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<14>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4109_1) );
	NAND2X1 NAND2X1_2574 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4108_1), .B(dp.rf._abc_6362_n4109_1), .Y(dp.rf._abc_6362_n3684) );
	NAND2X1 NAND2X1_2575 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4111_1) );
	NAND2X1 NAND2X1_2576 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<15>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4112_1) );
	NAND2X1 NAND2X1_2577 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4111_1), .B(dp.rf._abc_6362_n4112_1), .Y(dp.rf._abc_6362_n3685) );
	NAND2X1 NAND2X1_2578 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4114_1) );
	NAND2X1 NAND2X1_2579 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<16>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4115_1) );
	NAND2X1 NAND2X1_2580 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4114_1), .B(dp.rf._abc_6362_n4115_1), .Y(dp.rf._abc_6362_n3686) );
	NAND2X1 NAND2X1_2581 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4117_1) );
	NAND2X1 NAND2X1_2582 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<17>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4118_1) );
	NAND2X1 NAND2X1_2583 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4117_1), .B(dp.rf._abc_6362_n4118_1), .Y(dp.rf._abc_6362_n3687) );
	NAND2X1 NAND2X1_2584 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4120_1) );
	NAND2X1 NAND2X1_2585 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<18>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4121_1) );
	NAND2X1 NAND2X1_2586 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4120_1), .B(dp.rf._abc_6362_n4121_1), .Y(dp.rf._abc_6362_n3688) );
	NAND2X1 NAND2X1_2587 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4123_1) );
	NAND2X1 NAND2X1_2588 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<19>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4124_1) );
	NAND2X1 NAND2X1_2589 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4123_1), .B(dp.rf._abc_6362_n4124_1), .Y(dp.rf._abc_6362_n3689) );
	NAND2X1 NAND2X1_2590 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4126) );
	NAND2X1 NAND2X1_2591 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<20>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4127_1) );
	NAND2X1 NAND2X1_2592 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4126), .B(dp.rf._abc_6362_n4127_1), .Y(dp.rf._abc_6362_n3690) );
	NAND2X1 NAND2X1_2593 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4129_1) );
	NAND2X1 NAND2X1_2594 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<21>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4130) );
	NAND2X1 NAND2X1_2595 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4129_1), .B(dp.rf._abc_6362_n4130), .Y(dp.rf._abc_6362_n3691) );
	NAND2X1 NAND2X1_2596 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4132) );
	NAND2X1 NAND2X1_2597 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<22>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4133_1) );
	NAND2X1 NAND2X1_2598 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4132), .B(dp.rf._abc_6362_n4133_1), .Y(dp.rf._abc_6362_n3692) );
	NAND2X1 NAND2X1_2599 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4135_1) );
	NAND2X1 NAND2X1_2600 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<23>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4136) );
	NAND2X1 NAND2X1_2601 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4135_1), .B(dp.rf._abc_6362_n4136), .Y(dp.rf._abc_6362_n3693) );
	NAND2X1 NAND2X1_2602 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4138) );
	NAND2X1 NAND2X1_2603 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<24>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4139_1) );
	NAND2X1 NAND2X1_2604 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4138), .B(dp.rf._abc_6362_n4139_1), .Y(dp.rf._abc_6362_n3694) );
	NAND2X1 NAND2X1_2605 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4141_1) );
	NAND2X1 NAND2X1_2606 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<25>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4142) );
	NAND2X1 NAND2X1_2607 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4141_1), .B(dp.rf._abc_6362_n4142), .Y(dp.rf._abc_6362_n3695) );
	NAND2X1 NAND2X1_2608 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4144) );
	NAND2X1 NAND2X1_2609 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<26>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4145_1) );
	NAND2X1 NAND2X1_2610 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4144), .B(dp.rf._abc_6362_n4145_1), .Y(dp.rf._abc_6362_n3696) );
	NAND2X1 NAND2X1_2611 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4147_1) );
	NAND2X1 NAND2X1_2612 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<27>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4148) );
	NAND2X1 NAND2X1_2613 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4147_1), .B(dp.rf._abc_6362_n4148), .Y(dp.rf._abc_6362_n3697) );
	NAND2X1 NAND2X1_2614 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4150) );
	NAND2X1 NAND2X1_2615 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<28>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4151_1) );
	NAND2X1 NAND2X1_2616 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4150), .B(dp.rf._abc_6362_n4151_1), .Y(dp.rf._abc_6362_n3698) );
	NAND2X1 NAND2X1_2617 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4153_1) );
	NAND2X1 NAND2X1_2618 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<29>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4154) );
	NAND2X1 NAND2X1_2619 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4153_1), .B(dp.rf._abc_6362_n4154), .Y(dp.rf._abc_6362_n3699) );
	NAND2X1 NAND2X1_2620 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4156) );
	NAND2X1 NAND2X1_2621 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<30>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4157_1) );
	NAND2X1 NAND2X1_2622 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4156), .B(dp.rf._abc_6362_n4157_1), .Y(dp.rf._abc_6362_n3700) );
	NAND2X1 NAND2X1_2623 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n4064_1), .Y(dp.rf._abc_6362_n4159_1) );
	NAND2X1 NAND2X1_2624 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_27_<31>), .B(dp.rf._abc_6362_n4066_1), .Y(dp.rf._abc_6362_n4160) );
	NAND2X1 NAND2X1_2625 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4159_1), .B(dp.rf._abc_6362_n4160), .Y(dp.rf._abc_6362_n3701) );
	NOR2X1 NOR2X1_212 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n2477), .Y(dp.rf._abc_6362_n4162) );
	NAND2X1 NAND2X1_2626 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4163_1) );
	INVX8 INVX8_25 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4164) );
	NAND2X1 NAND2X1_2627 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<0>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4165_1) );
	NAND2X1 NAND2X1_2628 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4163_1), .B(dp.rf._abc_6362_n4165_1), .Y(dp.rf._abc_6362_n3702) );
	NAND2X1 NAND2X1_2629 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4167_1) );
	NAND2X1 NAND2X1_2630 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<1>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4168) );
	NAND2X1 NAND2X1_2631 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4167_1), .B(dp.rf._abc_6362_n4168), .Y(dp.rf._abc_6362_n3703) );
	NAND2X1 NAND2X1_2632 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4170) );
	NAND2X1 NAND2X1_2633 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<2>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4171_1) );
	NAND2X1 NAND2X1_2634 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4170), .B(dp.rf._abc_6362_n4171_1), .Y(dp.rf._abc_6362_n3704) );
	NAND2X1 NAND2X1_2635 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4173_1) );
	NAND2X1 NAND2X1_2636 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<3>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4174) );
	NAND2X1 NAND2X1_2637 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4173_1), .B(dp.rf._abc_6362_n4174), .Y(dp.rf._abc_6362_n3705) );
	NAND2X1 NAND2X1_2638 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4176) );
	NAND2X1 NAND2X1_2639 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<4>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4177_1) );
	NAND2X1 NAND2X1_2640 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4176), .B(dp.rf._abc_6362_n4177_1), .Y(dp.rf._abc_6362_n3706) );
	NAND2X1 NAND2X1_2641 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4179_1) );
	NAND2X1 NAND2X1_2642 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<5>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4180) );
	NAND2X1 NAND2X1_2643 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4179_1), .B(dp.rf._abc_6362_n4180), .Y(dp.rf._abc_6362_n3707) );
	NAND2X1 NAND2X1_2644 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4182) );
	NAND2X1 NAND2X1_2645 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<6>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4183_1) );
	NAND2X1 NAND2X1_2646 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4182), .B(dp.rf._abc_6362_n4183_1), .Y(dp.rf._abc_6362_n3708) );
	NAND2X1 NAND2X1_2647 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4185_1) );
	NAND2X1 NAND2X1_2648 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<7>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4186) );
	NAND2X1 NAND2X1_2649 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4185_1), .B(dp.rf._abc_6362_n4186), .Y(dp.rf._abc_6362_n3709) );
	NAND2X1 NAND2X1_2650 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4188) );
	NAND2X1 NAND2X1_2651 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<8>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4189_1) );
	NAND2X1 NAND2X1_2652 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4188), .B(dp.rf._abc_6362_n4189_1), .Y(dp.rf._abc_6362_n3710) );
	NAND2X1 NAND2X1_2653 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4191_1) );
	NAND2X1 NAND2X1_2654 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<9>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4192_1) );
	NAND2X1 NAND2X1_2655 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4191_1), .B(dp.rf._abc_6362_n4192_1), .Y(dp.rf._abc_6362_n3711) );
	NAND2X1 NAND2X1_2656 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4194_1) );
	NAND2X1 NAND2X1_2657 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<10>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4195_1) );
	NAND2X1 NAND2X1_2658 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4194_1), .B(dp.rf._abc_6362_n4195_1), .Y(dp.rf._abc_6362_n3712) );
	NAND2X1 NAND2X1_2659 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4197_1) );
	NAND2X1 NAND2X1_2660 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<11>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4198_1) );
	NAND2X1 NAND2X1_2661 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4197_1), .B(dp.rf._abc_6362_n4198_1), .Y(dp.rf._abc_6362_n3713) );
	NAND2X1 NAND2X1_2662 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4200_1) );
	NAND2X1 NAND2X1_2663 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<12>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4201_1) );
	NAND2X1 NAND2X1_2664 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4200_1), .B(dp.rf._abc_6362_n4201_1), .Y(dp.rf._abc_6362_n3714) );
	NAND2X1 NAND2X1_2665 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4203_1) );
	NAND2X1 NAND2X1_2666 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<13>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4204_1) );
	NAND2X1 NAND2X1_2667 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4203_1), .B(dp.rf._abc_6362_n4204_1), .Y(dp.rf._abc_6362_n3715) );
	NAND2X1 NAND2X1_2668 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4206_1) );
	NAND2X1 NAND2X1_2669 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<14>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4207_1) );
	NAND2X1 NAND2X1_2670 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4206_1), .B(dp.rf._abc_6362_n4207_1), .Y(dp.rf._abc_6362_n3716) );
	NAND2X1 NAND2X1_2671 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4209_1) );
	NAND2X1 NAND2X1_2672 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<15>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4210_1) );
	NAND2X1 NAND2X1_2673 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4209_1), .B(dp.rf._abc_6362_n4210_1), .Y(dp.rf._abc_6362_n3717) );
	NAND2X1 NAND2X1_2674 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4212_1) );
	NAND2X1 NAND2X1_2675 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<16>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4213_1) );
	NAND2X1 NAND2X1_2676 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4212_1), .B(dp.rf._abc_6362_n4213_1), .Y(dp.rf._abc_6362_n3718) );
	NAND2X1 NAND2X1_2677 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4215_1) );
	NAND2X1 NAND2X1_2678 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<17>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4216_1) );
	NAND2X1 NAND2X1_2679 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4215_1), .B(dp.rf._abc_6362_n4216_1), .Y(dp.rf._abc_6362_n3719) );
	NAND2X1 NAND2X1_2680 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4218_1) );
	NAND2X1 NAND2X1_2681 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<18>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4219_1) );
	NAND2X1 NAND2X1_2682 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4218_1), .B(dp.rf._abc_6362_n4219_1), .Y(dp.rf._abc_6362_n3720) );
	NAND2X1 NAND2X1_2683 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4221_1) );
	NAND2X1 NAND2X1_2684 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<19>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4222) );
	NAND2X1 NAND2X1_2685 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4221_1), .B(dp.rf._abc_6362_n4222), .Y(dp.rf._abc_6362_n3721) );
	NAND2X1 NAND2X1_2686 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4224) );
	NAND2X1 NAND2X1_2687 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<20>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4225) );
	NAND2X1 NAND2X1_2688 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4224), .B(dp.rf._abc_6362_n4225), .Y(dp.rf._abc_6362_n3722) );
	NAND2X1 NAND2X1_2689 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4227) );
	NAND2X1 NAND2X1_2690 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<21>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4228) );
	NAND2X1 NAND2X1_2691 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4227), .B(dp.rf._abc_6362_n4228), .Y(dp.rf._abc_6362_n3723) );
	NAND2X1 NAND2X1_2692 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4230) );
	NAND2X1 NAND2X1_2693 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<22>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4231) );
	NAND2X1 NAND2X1_2694 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4230), .B(dp.rf._abc_6362_n4231), .Y(dp.rf._abc_6362_n3724) );
	NAND2X1 NAND2X1_2695 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4233) );
	NAND2X1 NAND2X1_2696 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<23>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4234) );
	NAND2X1 NAND2X1_2697 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4233), .B(dp.rf._abc_6362_n4234), .Y(dp.rf._abc_6362_n3725) );
	NAND2X1 NAND2X1_2698 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4236) );
	NAND2X1 NAND2X1_2699 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<24>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4237) );
	NAND2X1 NAND2X1_2700 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4236), .B(dp.rf._abc_6362_n4237), .Y(dp.rf._abc_6362_n3726) );
	NAND2X1 NAND2X1_2701 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4239) );
	NAND2X1 NAND2X1_2702 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<25>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4240) );
	NAND2X1 NAND2X1_2703 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4239), .B(dp.rf._abc_6362_n4240), .Y(dp.rf._abc_6362_n3727) );
	NAND2X1 NAND2X1_2704 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4242) );
	NAND2X1 NAND2X1_2705 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<26>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4243) );
	NAND2X1 NAND2X1_2706 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4242), .B(dp.rf._abc_6362_n4243), .Y(dp.rf._abc_6362_n3728) );
	NAND2X1 NAND2X1_2707 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4245) );
	NAND2X1 NAND2X1_2708 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<27>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4246) );
	NAND2X1 NAND2X1_2709 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4245), .B(dp.rf._abc_6362_n4246), .Y(dp.rf._abc_6362_n3729) );
	NAND2X1 NAND2X1_2710 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4248) );
	NAND2X1 NAND2X1_2711 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<28>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4249) );
	NAND2X1 NAND2X1_2712 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4248), .B(dp.rf._abc_6362_n4249), .Y(dp.rf._abc_6362_n3730) );
	NAND2X1 NAND2X1_2713 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4251) );
	NAND2X1 NAND2X1_2714 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<29>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4252) );
	NAND2X1 NAND2X1_2715 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4251), .B(dp.rf._abc_6362_n4252), .Y(dp.rf._abc_6362_n3731) );
	NAND2X1 NAND2X1_2716 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4254) );
	NAND2X1 NAND2X1_2717 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<30>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4255) );
	NAND2X1 NAND2X1_2718 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4254), .B(dp.rf._abc_6362_n4255), .Y(dp.rf._abc_6362_n3732) );
	NAND2X1 NAND2X1_2719 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n4162), .Y(dp.rf._abc_6362_n4257) );
	NAND2X1 NAND2X1_2720 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<31>), .B(dp.rf._abc_6362_n4164), .Y(dp.rf._abc_6362_n4258) );
	NAND2X1 NAND2X1_2721 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4257), .B(dp.rf._abc_6362_n4258), .Y(dp.rf._abc_6362_n3733) );
	NOR2X1 NOR2X1_213 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n2577), .Y(dp.rf._abc_6362_n4260) );
	NAND2X1 NAND2X1_2722 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4261) );
	INVX8 INVX8_26 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4262) );
	NAND2X1 NAND2X1_2723 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<0>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4263) );
	NAND2X1 NAND2X1_2724 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4261), .B(dp.rf._abc_6362_n4263), .Y(dp.rf._abc_6362_n3734) );
	NAND2X1 NAND2X1_2725 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4265) );
	NAND2X1 NAND2X1_2726 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<1>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4266) );
	NAND2X1 NAND2X1_2727 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4265), .B(dp.rf._abc_6362_n4266), .Y(dp.rf._abc_6362_n3735) );
	NAND2X1 NAND2X1_2728 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4268) );
	NAND2X1 NAND2X1_2729 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<2>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4269) );
	NAND2X1 NAND2X1_2730 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4268), .B(dp.rf._abc_6362_n4269), .Y(dp.rf._abc_6362_n3736) );
	NAND2X1 NAND2X1_2731 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4271) );
	NAND2X1 NAND2X1_2732 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<3>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4272) );
	NAND2X1 NAND2X1_2733 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4271), .B(dp.rf._abc_6362_n4272), .Y(dp.rf._abc_6362_n3737) );
	NAND2X1 NAND2X1_2734 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4274) );
	NAND2X1 NAND2X1_2735 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<4>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4275) );
	NAND2X1 NAND2X1_2736 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4274), .B(dp.rf._abc_6362_n4275), .Y(dp.rf._abc_6362_n3738) );
	NAND2X1 NAND2X1_2737 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4277) );
	NAND2X1 NAND2X1_2738 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<5>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4278) );
	NAND2X1 NAND2X1_2739 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4277), .B(dp.rf._abc_6362_n4278), .Y(dp.rf._abc_6362_n3739) );
	NAND2X1 NAND2X1_2740 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4280) );
	NAND2X1 NAND2X1_2741 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<6>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4281) );
	NAND2X1 NAND2X1_2742 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4280), .B(dp.rf._abc_6362_n4281), .Y(dp.rf._abc_6362_n3740) );
	NAND2X1 NAND2X1_2743 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4283) );
	NAND2X1 NAND2X1_2744 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<7>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4284) );
	NAND2X1 NAND2X1_2745 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4283), .B(dp.rf._abc_6362_n4284), .Y(dp.rf._abc_6362_n3741) );
	NAND2X1 NAND2X1_2746 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4286) );
	NAND2X1 NAND2X1_2747 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<8>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4287) );
	NAND2X1 NAND2X1_2748 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4286), .B(dp.rf._abc_6362_n4287), .Y(dp.rf._abc_6362_n3742) );
	NAND2X1 NAND2X1_2749 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4289) );
	NAND2X1 NAND2X1_2750 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<9>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4290) );
	NAND2X1 NAND2X1_2751 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4289), .B(dp.rf._abc_6362_n4290), .Y(dp.rf._abc_6362_n3743) );
	NAND2X1 NAND2X1_2752 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4292) );
	NAND2X1 NAND2X1_2753 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<10>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4293) );
	NAND2X1 NAND2X1_2754 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4292), .B(dp.rf._abc_6362_n4293), .Y(dp.rf._abc_6362_n3744) );
	NAND2X1 NAND2X1_2755 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4295) );
	NAND2X1 NAND2X1_2756 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<11>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4296) );
	NAND2X1 NAND2X1_2757 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4295), .B(dp.rf._abc_6362_n4296), .Y(dp.rf._abc_6362_n3745) );
	NAND2X1 NAND2X1_2758 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4298) );
	NAND2X1 NAND2X1_2759 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<12>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4299) );
	NAND2X1 NAND2X1_2760 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4298), .B(dp.rf._abc_6362_n4299), .Y(dp.rf._abc_6362_n3746) );
	NAND2X1 NAND2X1_2761 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4301) );
	NAND2X1 NAND2X1_2762 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<13>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4302) );
	NAND2X1 NAND2X1_2763 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4301), .B(dp.rf._abc_6362_n4302), .Y(dp.rf._abc_6362_n3747) );
	NAND2X1 NAND2X1_2764 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4304) );
	NAND2X1 NAND2X1_2765 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<14>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4305) );
	NAND2X1 NAND2X1_2766 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4304), .B(dp.rf._abc_6362_n4305), .Y(dp.rf._abc_6362_n3748) );
	NAND2X1 NAND2X1_2767 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4307) );
	NAND2X1 NAND2X1_2768 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<15>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4308) );
	NAND2X1 NAND2X1_2769 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4307), .B(dp.rf._abc_6362_n4308), .Y(dp.rf._abc_6362_n3749) );
	NAND2X1 NAND2X1_2770 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4310) );
	NAND2X1 NAND2X1_2771 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<16>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4311) );
	NAND2X1 NAND2X1_2772 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4310), .B(dp.rf._abc_6362_n4311), .Y(dp.rf._abc_6362_n3750) );
	NAND2X1 NAND2X1_2773 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4313) );
	NAND2X1 NAND2X1_2774 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<17>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4314) );
	NAND2X1 NAND2X1_2775 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4313), .B(dp.rf._abc_6362_n4314), .Y(dp.rf._abc_6362_n3751) );
	NAND2X1 NAND2X1_2776 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4316) );
	NAND2X1 NAND2X1_2777 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<18>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4317) );
	NAND2X1 NAND2X1_2778 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4316), .B(dp.rf._abc_6362_n4317), .Y(dp.rf._abc_6362_n3752) );
	NAND2X1 NAND2X1_2779 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4319) );
	NAND2X1 NAND2X1_2780 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<19>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4320) );
	NAND2X1 NAND2X1_2781 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4319), .B(dp.rf._abc_6362_n4320), .Y(dp.rf._abc_6362_n3753) );
	NAND2X1 NAND2X1_2782 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4322) );
	NAND2X1 NAND2X1_2783 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<20>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4323) );
	NAND2X1 NAND2X1_2784 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4322), .B(dp.rf._abc_6362_n4323), .Y(dp.rf._abc_6362_n3754) );
	NAND2X1 NAND2X1_2785 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4325) );
	NAND2X1 NAND2X1_2786 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<21>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4326) );
	NAND2X1 NAND2X1_2787 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4325), .B(dp.rf._abc_6362_n4326), .Y(dp.rf._abc_6362_n3755) );
	NAND2X1 NAND2X1_2788 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4328) );
	NAND2X1 NAND2X1_2789 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<22>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4329) );
	NAND2X1 NAND2X1_2790 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4328), .B(dp.rf._abc_6362_n4329), .Y(dp.rf._abc_6362_n3756) );
	NAND2X1 NAND2X1_2791 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4331) );
	NAND2X1 NAND2X1_2792 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<23>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4332) );
	NAND2X1 NAND2X1_2793 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4331), .B(dp.rf._abc_6362_n4332), .Y(dp.rf._abc_6362_n3757) );
	NAND2X1 NAND2X1_2794 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4334) );
	NAND2X1 NAND2X1_2795 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<24>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4335) );
	NAND2X1 NAND2X1_2796 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4334), .B(dp.rf._abc_6362_n4335), .Y(dp.rf._abc_6362_n3758) );
	NAND2X1 NAND2X1_2797 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4337) );
	NAND2X1 NAND2X1_2798 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<25>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4338) );
	NAND2X1 NAND2X1_2799 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4337), .B(dp.rf._abc_6362_n4338), .Y(dp.rf._abc_6362_n3759) );
	NAND2X1 NAND2X1_2800 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4340) );
	NAND2X1 NAND2X1_2801 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<26>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4341) );
	NAND2X1 NAND2X1_2802 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4340), .B(dp.rf._abc_6362_n4341), .Y(dp.rf._abc_6362_n3760) );
	NAND2X1 NAND2X1_2803 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4343) );
	NAND2X1 NAND2X1_2804 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<27>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4344) );
	NAND2X1 NAND2X1_2805 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4343), .B(dp.rf._abc_6362_n4344), .Y(dp.rf._abc_6362_n3761) );
	NAND2X1 NAND2X1_2806 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4346) );
	NAND2X1 NAND2X1_2807 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<28>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4347) );
	NAND2X1 NAND2X1_2808 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4346), .B(dp.rf._abc_6362_n4347), .Y(dp.rf._abc_6362_n3762) );
	NAND2X1 NAND2X1_2809 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4349) );
	NAND2X1 NAND2X1_2810 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<29>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4350) );
	NAND2X1 NAND2X1_2811 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4349), .B(dp.rf._abc_6362_n4350), .Y(dp.rf._abc_6362_n3763) );
	NAND2X1 NAND2X1_2812 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4352) );
	NAND2X1 NAND2X1_2813 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<30>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4353) );
	NAND2X1 NAND2X1_2814 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4352), .B(dp.rf._abc_6362_n4353), .Y(dp.rf._abc_6362_n3764) );
	NAND2X1 NAND2X1_2815 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n4260), .Y(dp.rf._abc_6362_n4355) );
	NAND2X1 NAND2X1_2816 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_29_<31>), .B(dp.rf._abc_6362_n4262), .Y(dp.rf._abc_6362_n4356) );
	NAND2X1 NAND2X1_2817 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4355), .B(dp.rf._abc_6362_n4356), .Y(dp.rf._abc_6362_n3765) );
	NOR2X1 NOR2X1_214 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n3073_1), .Y(dp.rf._abc_6362_n4358) );
	NAND2X1 NAND2X1_2818 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4359) );
	INVX8 INVX8_27 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4360) );
	NAND2X1 NAND2X1_2819 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<0>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4361) );
	NAND2X1 NAND2X1_2820 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4359), .B(dp.rf._abc_6362_n4361), .Y(dp.rf._abc_6362_n3766) );
	NAND2X1 NAND2X1_2821 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4363) );
	NAND2X1 NAND2X1_2822 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<1>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4364) );
	NAND2X1 NAND2X1_2823 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4363), .B(dp.rf._abc_6362_n4364), .Y(dp.rf._abc_6362_n3767) );
	NAND2X1 NAND2X1_2824 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4366) );
	NAND2X1 NAND2X1_2825 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<2>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4367) );
	NAND2X1 NAND2X1_2826 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4366), .B(dp.rf._abc_6362_n4367), .Y(dp.rf._abc_6362_n3768) );
	NAND2X1 NAND2X1_2827 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4369) );
	NAND2X1 NAND2X1_2828 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<3>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4370) );
	NAND2X1 NAND2X1_2829 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4369), .B(dp.rf._abc_6362_n4370), .Y(dp.rf._abc_6362_n3769) );
	NAND2X1 NAND2X1_2830 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4372) );
	NAND2X1 NAND2X1_2831 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<4>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4373) );
	NAND2X1 NAND2X1_2832 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4372), .B(dp.rf._abc_6362_n4373), .Y(dp.rf._abc_6362_n3770) );
	NAND2X1 NAND2X1_2833 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4375) );
	NAND2X1 NAND2X1_2834 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<5>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4376) );
	NAND2X1 NAND2X1_2835 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4375), .B(dp.rf._abc_6362_n4376), .Y(dp.rf._abc_6362_n3771) );
	NAND2X1 NAND2X1_2836 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4378) );
	NAND2X1 NAND2X1_2837 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<6>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4379) );
	NAND2X1 NAND2X1_2838 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4378), .B(dp.rf._abc_6362_n4379), .Y(dp.rf._abc_6362_n3772) );
	NAND2X1 NAND2X1_2839 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4381) );
	NAND2X1 NAND2X1_2840 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<7>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4382) );
	NAND2X1 NAND2X1_2841 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4381), .B(dp.rf._abc_6362_n4382), .Y(dp.rf._abc_6362_n3773) );
	NAND2X1 NAND2X1_2842 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4384) );
	NAND2X1 NAND2X1_2843 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<8>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4385) );
	NAND2X1 NAND2X1_2844 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4384), .B(dp.rf._abc_6362_n4385), .Y(dp.rf._abc_6362_n3774) );
	NAND2X1 NAND2X1_2845 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4387) );
	NAND2X1 NAND2X1_2846 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<9>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4388) );
	NAND2X1 NAND2X1_2847 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4387), .B(dp.rf._abc_6362_n4388), .Y(dp.rf._abc_6362_n3775) );
	NAND2X1 NAND2X1_2848 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4390) );
	NAND2X1 NAND2X1_2849 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<10>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4391) );
	NAND2X1 NAND2X1_2850 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4390), .B(dp.rf._abc_6362_n4391), .Y(dp.rf._abc_6362_n3776) );
	NAND2X1 NAND2X1_2851 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4393) );
	NAND2X1 NAND2X1_2852 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<11>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4394) );
	NAND2X1 NAND2X1_2853 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4393), .B(dp.rf._abc_6362_n4394), .Y(dp.rf._abc_6362_n3777) );
	NAND2X1 NAND2X1_2854 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4396) );
	NAND2X1 NAND2X1_2855 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<12>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4397) );
	NAND2X1 NAND2X1_2856 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4396), .B(dp.rf._abc_6362_n4397), .Y(dp.rf._abc_6362_n3778) );
	NAND2X1 NAND2X1_2857 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4399) );
	NAND2X1 NAND2X1_2858 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<13>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4400) );
	NAND2X1 NAND2X1_2859 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4399), .B(dp.rf._abc_6362_n4400), .Y(dp.rf._abc_6362_n3779) );
	NAND2X1 NAND2X1_2860 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4402) );
	NAND2X1 NAND2X1_2861 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<14>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4403) );
	NAND2X1 NAND2X1_2862 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4402), .B(dp.rf._abc_6362_n4403), .Y(dp.rf._abc_6362_n3780) );
	NAND2X1 NAND2X1_2863 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4405) );
	NAND2X1 NAND2X1_2864 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<15>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4406) );
	NAND2X1 NAND2X1_2865 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4405), .B(dp.rf._abc_6362_n4406), .Y(dp.rf._abc_6362_n3781) );
	NAND2X1 NAND2X1_2866 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4408) );
	NAND2X1 NAND2X1_2867 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<16>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4409) );
	NAND2X1 NAND2X1_2868 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4408), .B(dp.rf._abc_6362_n4409), .Y(dp.rf._abc_6362_n3782) );
	NAND2X1 NAND2X1_2869 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4411) );
	NAND2X1 NAND2X1_2870 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<17>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4412) );
	NAND2X1 NAND2X1_2871 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4411), .B(dp.rf._abc_6362_n4412), .Y(dp.rf._abc_6362_n3783) );
	NAND2X1 NAND2X1_2872 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4414) );
	NAND2X1 NAND2X1_2873 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<18>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4415) );
	NAND2X1 NAND2X1_2874 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4414), .B(dp.rf._abc_6362_n4415), .Y(dp.rf._abc_6362_n3784) );
	NAND2X1 NAND2X1_2875 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4417) );
	NAND2X1 NAND2X1_2876 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<19>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4418) );
	NAND2X1 NAND2X1_2877 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4417), .B(dp.rf._abc_6362_n4418), .Y(dp.rf._abc_6362_n3785) );
	NAND2X1 NAND2X1_2878 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4420) );
	NAND2X1 NAND2X1_2879 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<20>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4421) );
	NAND2X1 NAND2X1_2880 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4420), .B(dp.rf._abc_6362_n4421), .Y(dp.rf._abc_6362_n3786) );
	NAND2X1 NAND2X1_2881 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4423) );
	NAND2X1 NAND2X1_2882 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<21>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4424) );
	NAND2X1 NAND2X1_2883 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4423), .B(dp.rf._abc_6362_n4424), .Y(dp.rf._abc_6362_n3787) );
	NAND2X1 NAND2X1_2884 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4426) );
	NAND2X1 NAND2X1_2885 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<22>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4427) );
	NAND2X1 NAND2X1_2886 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4426), .B(dp.rf._abc_6362_n4427), .Y(dp.rf._abc_6362_n3788) );
	NAND2X1 NAND2X1_2887 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4429) );
	NAND2X1 NAND2X1_2888 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<23>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4430) );
	NAND2X1 NAND2X1_2889 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4429), .B(dp.rf._abc_6362_n4430), .Y(dp.rf._abc_6362_n3789) );
	NAND2X1 NAND2X1_2890 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4432) );
	NAND2X1 NAND2X1_2891 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<24>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4433) );
	NAND2X1 NAND2X1_2892 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4432), .B(dp.rf._abc_6362_n4433), .Y(dp.rf._abc_6362_n3790) );
	NAND2X1 NAND2X1_2893 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4435) );
	NAND2X1 NAND2X1_2894 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<25>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4436) );
	NAND2X1 NAND2X1_2895 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4435), .B(dp.rf._abc_6362_n4436), .Y(dp.rf._abc_6362_n3791) );
	NAND2X1 NAND2X1_2896 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4438) );
	NAND2X1 NAND2X1_2897 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<26>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4439) );
	NAND2X1 NAND2X1_2898 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4438), .B(dp.rf._abc_6362_n4439), .Y(dp.rf._abc_6362_n3792) );
	NAND2X1 NAND2X1_2899 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4441) );
	NAND2X1 NAND2X1_2900 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<27>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4442) );
	NAND2X1 NAND2X1_2901 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4441), .B(dp.rf._abc_6362_n4442), .Y(dp.rf._abc_6362_n3793) );
	NAND2X1 NAND2X1_2902 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4444) );
	NAND2X1 NAND2X1_2903 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<28>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4445) );
	NAND2X1 NAND2X1_2904 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4444), .B(dp.rf._abc_6362_n4445), .Y(dp.rf._abc_6362_n3794) );
	NAND2X1 NAND2X1_2905 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4447) );
	NAND2X1 NAND2X1_2906 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<29>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4448) );
	NAND2X1 NAND2X1_2907 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4447), .B(dp.rf._abc_6362_n4448), .Y(dp.rf._abc_6362_n3795) );
	NAND2X1 NAND2X1_2908 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4450) );
	NAND2X1 NAND2X1_2909 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<30>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4451) );
	NAND2X1 NAND2X1_2910 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4450), .B(dp.rf._abc_6362_n4451), .Y(dp.rf._abc_6362_n3796) );
	NAND2X1 NAND2X1_2911 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n4358), .Y(dp.rf._abc_6362_n4453) );
	NAND2X1 NAND2X1_2912 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<31>), .B(dp.rf._abc_6362_n4360), .Y(dp.rf._abc_6362_n4454) );
	NAND2X1 NAND2X1_2913 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4453), .B(dp.rf._abc_6362_n4454), .Y(dp.rf._abc_6362_n3797) );
	NOR2X1 NOR2X1_215 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n2676), .Y(dp.rf._abc_6362_n4456) );
	NAND2X1 NAND2X1_2914 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4457) );
	INVX8 INVX8_28 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4458) );
	NAND2X1 NAND2X1_2915 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<0>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4459) );
	NAND2X1 NAND2X1_2916 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4457), .B(dp.rf._abc_6362_n4459), .Y(dp.rf._abc_6362_n3798) );
	NAND2X1 NAND2X1_2917 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4461) );
	NAND2X1 NAND2X1_2918 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<1>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4462) );
	NAND2X1 NAND2X1_2919 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4461), .B(dp.rf._abc_6362_n4462), .Y(dp.rf._abc_6362_n3799) );
	NAND2X1 NAND2X1_2920 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4464) );
	NAND2X1 NAND2X1_2921 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<2>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4465) );
	NAND2X1 NAND2X1_2922 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4464), .B(dp.rf._abc_6362_n4465), .Y(dp.rf._abc_6362_n3800) );
	NAND2X1 NAND2X1_2923 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4467) );
	NAND2X1 NAND2X1_2924 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<3>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4468) );
	NAND2X1 NAND2X1_2925 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4467), .B(dp.rf._abc_6362_n4468), .Y(dp.rf._abc_6362_n3801) );
	NAND2X1 NAND2X1_2926 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4470) );
	NAND2X1 NAND2X1_2927 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<4>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4471) );
	NAND2X1 NAND2X1_2928 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4470), .B(dp.rf._abc_6362_n4471), .Y(dp.rf._abc_6362_n3802) );
	NAND2X1 NAND2X1_2929 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4473) );
	NAND2X1 NAND2X1_2930 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<5>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4474) );
	NAND2X1 NAND2X1_2931 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4473), .B(dp.rf._abc_6362_n4474), .Y(dp.rf._abc_6362_n3803) );
	NAND2X1 NAND2X1_2932 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4476) );
	NAND2X1 NAND2X1_2933 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<6>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4477) );
	NAND2X1 NAND2X1_2934 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4476), .B(dp.rf._abc_6362_n4477), .Y(dp.rf._abc_6362_n3804) );
	NAND2X1 NAND2X1_2935 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4479) );
	NAND2X1 NAND2X1_2936 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<7>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4480) );
	NAND2X1 NAND2X1_2937 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4479), .B(dp.rf._abc_6362_n4480), .Y(dp.rf._abc_6362_n3805) );
	NAND2X1 NAND2X1_2938 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4482) );
	NAND2X1 NAND2X1_2939 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<8>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4483) );
	NAND2X1 NAND2X1_2940 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4482), .B(dp.rf._abc_6362_n4483), .Y(dp.rf._abc_6362_n3806) );
	NAND2X1 NAND2X1_2941 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4485) );
	NAND2X1 NAND2X1_2942 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<9>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4486) );
	NAND2X1 NAND2X1_2943 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4485), .B(dp.rf._abc_6362_n4486), .Y(dp.rf._abc_6362_n3807) );
	NAND2X1 NAND2X1_2944 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4488) );
	NAND2X1 NAND2X1_2945 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<10>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4489) );
	NAND2X1 NAND2X1_2946 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4488), .B(dp.rf._abc_6362_n4489), .Y(dp.rf._abc_6362_n3808) );
	NAND2X1 NAND2X1_2947 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4491) );
	NAND2X1 NAND2X1_2948 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<11>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4492) );
	NAND2X1 NAND2X1_2949 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4491), .B(dp.rf._abc_6362_n4492), .Y(dp.rf._abc_6362_n3809) );
	NAND2X1 NAND2X1_2950 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4494) );
	NAND2X1 NAND2X1_2951 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<12>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4495) );
	NAND2X1 NAND2X1_2952 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4494), .B(dp.rf._abc_6362_n4495), .Y(dp.rf._abc_6362_n3810) );
	NAND2X1 NAND2X1_2953 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4497) );
	NAND2X1 NAND2X1_2954 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<13>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4498) );
	NAND2X1 NAND2X1_2955 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4497), .B(dp.rf._abc_6362_n4498), .Y(dp.rf._abc_6362_n3811) );
	NAND2X1 NAND2X1_2956 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4500) );
	NAND2X1 NAND2X1_2957 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<14>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4501) );
	NAND2X1 NAND2X1_2958 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4500), .B(dp.rf._abc_6362_n4501), .Y(dp.rf._abc_6362_n3812) );
	NAND2X1 NAND2X1_2959 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4503) );
	NAND2X1 NAND2X1_2960 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<15>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4504) );
	NAND2X1 NAND2X1_2961 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4503), .B(dp.rf._abc_6362_n4504), .Y(dp.rf._abc_6362_n3813) );
	NAND2X1 NAND2X1_2962 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4506) );
	NAND2X1 NAND2X1_2963 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<16>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4507) );
	NAND2X1 NAND2X1_2964 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4506), .B(dp.rf._abc_6362_n4507), .Y(dp.rf._abc_6362_n3814) );
	NAND2X1 NAND2X1_2965 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4509) );
	NAND2X1 NAND2X1_2966 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<17>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4510) );
	NAND2X1 NAND2X1_2967 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4509), .B(dp.rf._abc_6362_n4510), .Y(dp.rf._abc_6362_n3815) );
	NAND2X1 NAND2X1_2968 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4512) );
	NAND2X1 NAND2X1_2969 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<18>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4513) );
	NAND2X1 NAND2X1_2970 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4512), .B(dp.rf._abc_6362_n4513), .Y(dp.rf._abc_6362_n3816) );
	NAND2X1 NAND2X1_2971 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4515) );
	NAND2X1 NAND2X1_2972 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<19>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4516) );
	NAND2X1 NAND2X1_2973 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4515), .B(dp.rf._abc_6362_n4516), .Y(dp.rf._abc_6362_n3817) );
	NAND2X1 NAND2X1_2974 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4518) );
	NAND2X1 NAND2X1_2975 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<20>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4519) );
	NAND2X1 NAND2X1_2976 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4518), .B(dp.rf._abc_6362_n4519), .Y(dp.rf._abc_6362_n3818) );
	NAND2X1 NAND2X1_2977 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4521) );
	NAND2X1 NAND2X1_2978 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<21>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4522) );
	NAND2X1 NAND2X1_2979 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4521), .B(dp.rf._abc_6362_n4522), .Y(dp.rf._abc_6362_n3819) );
	NAND2X1 NAND2X1_2980 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4524) );
	NAND2X1 NAND2X1_2981 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<22>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4525) );
	NAND2X1 NAND2X1_2982 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4524), .B(dp.rf._abc_6362_n4525), .Y(dp.rf._abc_6362_n3820) );
	NAND2X1 NAND2X1_2983 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4527) );
	NAND2X1 NAND2X1_2984 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<23>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4528) );
	NAND2X1 NAND2X1_2985 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4527), .B(dp.rf._abc_6362_n4528), .Y(dp.rf._abc_6362_n3821) );
	NAND2X1 NAND2X1_2986 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4530) );
	NAND2X1 NAND2X1_2987 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<24>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4531) );
	NAND2X1 NAND2X1_2988 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4530), .B(dp.rf._abc_6362_n4531), .Y(dp.rf._abc_6362_n3822) );
	NAND2X1 NAND2X1_2989 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4533) );
	NAND2X1 NAND2X1_2990 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<25>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4534) );
	NAND2X1 NAND2X1_2991 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4533), .B(dp.rf._abc_6362_n4534), .Y(dp.rf._abc_6362_n3823) );
	NAND2X1 NAND2X1_2992 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4536) );
	NAND2X1 NAND2X1_2993 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<26>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4537) );
	NAND2X1 NAND2X1_2994 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4536), .B(dp.rf._abc_6362_n4537), .Y(dp.rf._abc_6362_n3824) );
	NAND2X1 NAND2X1_2995 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4539) );
	NAND2X1 NAND2X1_2996 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<27>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4540) );
	NAND2X1 NAND2X1_2997 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4539), .B(dp.rf._abc_6362_n4540), .Y(dp.rf._abc_6362_n3825) );
	NAND2X1 NAND2X1_2998 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4542) );
	NAND2X1 NAND2X1_2999 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<28>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4543) );
	NAND2X1 NAND2X1_3000 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4542), .B(dp.rf._abc_6362_n4543), .Y(dp.rf._abc_6362_n3826) );
	NAND2X1 NAND2X1_3001 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4545) );
	NAND2X1 NAND2X1_3002 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<29>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4546) );
	NAND2X1 NAND2X1_3003 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4545), .B(dp.rf._abc_6362_n4546), .Y(dp.rf._abc_6362_n3827) );
	NAND2X1 NAND2X1_3004 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4548) );
	NAND2X1 NAND2X1_3005 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<30>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4549) );
	NAND2X1 NAND2X1_3006 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4548), .B(dp.rf._abc_6362_n4549), .Y(dp.rf._abc_6362_n3828) );
	NAND2X1 NAND2X1_3007 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n4456), .Y(dp.rf._abc_6362_n4551) );
	NAND2X1 NAND2X1_3008 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<31>), .B(dp.rf._abc_6362_n4458), .Y(dp.rf._abc_6362_n4552) );
	NAND2X1 NAND2X1_3009 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4551), .B(dp.rf._abc_6362_n4552), .Y(dp.rf._abc_6362_n3829) );
	NOR2X1 NOR2X1_216 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2875), .B(dp.rf._abc_6362_n2775), .Y(dp.rf._abc_6362_n4554) );
	NAND2X1 NAND2X1_3010 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4555) );
	INVX8 INVX8_29 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4556) );
	NAND2X1 NAND2X1_3011 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<0>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4557) );
	NAND2X1 NAND2X1_3012 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4555), .B(dp.rf._abc_6362_n4557), .Y(dp.rf._abc_6362_n3830) );
	NAND2X1 NAND2X1_3013 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4559) );
	NAND2X1 NAND2X1_3014 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<1>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4560) );
	NAND2X1 NAND2X1_3015 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4559), .B(dp.rf._abc_6362_n4560), .Y(dp.rf._abc_6362_n3831) );
	NAND2X1 NAND2X1_3016 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4562) );
	NAND2X1 NAND2X1_3017 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<2>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4563) );
	NAND2X1 NAND2X1_3018 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4562), .B(dp.rf._abc_6362_n4563), .Y(dp.rf._abc_6362_n3832) );
	NAND2X1 NAND2X1_3019 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4565) );
	NAND2X1 NAND2X1_3020 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<3>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4566) );
	NAND2X1 NAND2X1_3021 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4565), .B(dp.rf._abc_6362_n4566), .Y(dp.rf._abc_6362_n3833) );
	NAND2X1 NAND2X1_3022 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4568) );
	NAND2X1 NAND2X1_3023 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<4>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4569) );
	NAND2X1 NAND2X1_3024 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4568), .B(dp.rf._abc_6362_n4569), .Y(dp.rf._abc_6362_n3834) );
	NAND2X1 NAND2X1_3025 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4571) );
	NAND2X1 NAND2X1_3026 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<5>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4572) );
	NAND2X1 NAND2X1_3027 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4571), .B(dp.rf._abc_6362_n4572), .Y(dp.rf._abc_6362_n3835) );
	NAND2X1 NAND2X1_3028 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4574) );
	NAND2X1 NAND2X1_3029 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<6>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4575) );
	NAND2X1 NAND2X1_3030 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4574), .B(dp.rf._abc_6362_n4575), .Y(dp.rf._abc_6362_n3836) );
	NAND2X1 NAND2X1_3031 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4577) );
	NAND2X1 NAND2X1_3032 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<7>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4578) );
	NAND2X1 NAND2X1_3033 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4577), .B(dp.rf._abc_6362_n4578), .Y(dp.rf._abc_6362_n3837) );
	NAND2X1 NAND2X1_3034 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4580) );
	NAND2X1 NAND2X1_3035 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<8>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4581) );
	NAND2X1 NAND2X1_3036 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4580), .B(dp.rf._abc_6362_n4581), .Y(dp.rf._abc_6362_n3838) );
	NAND2X1 NAND2X1_3037 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4583) );
	NAND2X1 NAND2X1_3038 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<9>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4584) );
	NAND2X1 NAND2X1_3039 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4583), .B(dp.rf._abc_6362_n4584), .Y(dp.rf._abc_6362_n3839) );
	NAND2X1 NAND2X1_3040 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4586) );
	NAND2X1 NAND2X1_3041 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<10>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4587) );
	NAND2X1 NAND2X1_3042 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4586), .B(dp.rf._abc_6362_n4587), .Y(dp.rf._abc_6362_n3840) );
	NAND2X1 NAND2X1_3043 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4589) );
	NAND2X1 NAND2X1_3044 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<11>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4590) );
	NAND2X1 NAND2X1_3045 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4589), .B(dp.rf._abc_6362_n4590), .Y(dp.rf._abc_6362_n3841) );
	NAND2X1 NAND2X1_3046 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4592) );
	NAND2X1 NAND2X1_3047 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<12>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4593) );
	NAND2X1 NAND2X1_3048 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4592), .B(dp.rf._abc_6362_n4593), .Y(dp.rf._abc_6362_n3842) );
	NAND2X1 NAND2X1_3049 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4595) );
	NAND2X1 NAND2X1_3050 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<13>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4596) );
	NAND2X1 NAND2X1_3051 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4595), .B(dp.rf._abc_6362_n4596), .Y(dp.rf._abc_6362_n3843) );
	NAND2X1 NAND2X1_3052 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4598) );
	NAND2X1 NAND2X1_3053 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<14>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4599) );
	NAND2X1 NAND2X1_3054 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4598), .B(dp.rf._abc_6362_n4599), .Y(dp.rf._abc_6362_n3844) );
	NAND2X1 NAND2X1_3055 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4601) );
	NAND2X1 NAND2X1_3056 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<15>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4602) );
	NAND2X1 NAND2X1_3057 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4601), .B(dp.rf._abc_6362_n4602), .Y(dp.rf._abc_6362_n3845) );
	NAND2X1 NAND2X1_3058 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4604) );
	NAND2X1 NAND2X1_3059 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<16>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4605) );
	NAND2X1 NAND2X1_3060 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4604), .B(dp.rf._abc_6362_n4605), .Y(dp.rf._abc_6362_n3846) );
	NAND2X1 NAND2X1_3061 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4607) );
	NAND2X1 NAND2X1_3062 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<17>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4608) );
	NAND2X1 NAND2X1_3063 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4607), .B(dp.rf._abc_6362_n4608), .Y(dp.rf._abc_6362_n3847) );
	NAND2X1 NAND2X1_3064 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4610) );
	NAND2X1 NAND2X1_3065 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<18>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4611) );
	NAND2X1 NAND2X1_3066 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4610), .B(dp.rf._abc_6362_n4611), .Y(dp.rf._abc_6362_n3848) );
	NAND2X1 NAND2X1_3067 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4613) );
	NAND2X1 NAND2X1_3068 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<19>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4614) );
	NAND2X1 NAND2X1_3069 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4613), .B(dp.rf._abc_6362_n4614), .Y(dp.rf._abc_6362_n3849) );
	NAND2X1 NAND2X1_3070 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4616) );
	NAND2X1 NAND2X1_3071 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<20>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4617) );
	NAND2X1 NAND2X1_3072 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4616), .B(dp.rf._abc_6362_n4617), .Y(dp.rf._abc_6362_n3850) );
	NAND2X1 NAND2X1_3073 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4619) );
	NAND2X1 NAND2X1_3074 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<21>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4620) );
	NAND2X1 NAND2X1_3075 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4619), .B(dp.rf._abc_6362_n4620), .Y(dp.rf._abc_6362_n3851) );
	NAND2X1 NAND2X1_3076 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4622) );
	NAND2X1 NAND2X1_3077 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<22>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4623) );
	NAND2X1 NAND2X1_3078 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4622), .B(dp.rf._abc_6362_n4623), .Y(dp.rf._abc_6362_n3852) );
	NAND2X1 NAND2X1_3079 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4625) );
	NAND2X1 NAND2X1_3080 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<23>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4626) );
	NAND2X1 NAND2X1_3081 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4625), .B(dp.rf._abc_6362_n4626), .Y(dp.rf._abc_6362_n3853) );
	NAND2X1 NAND2X1_3082 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4628) );
	NAND2X1 NAND2X1_3083 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<24>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4629) );
	NAND2X1 NAND2X1_3084 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4628), .B(dp.rf._abc_6362_n4629), .Y(dp.rf._abc_6362_n3854) );
	NAND2X1 NAND2X1_3085 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4631) );
	NAND2X1 NAND2X1_3086 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<25>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4632) );
	NAND2X1 NAND2X1_3087 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4631), .B(dp.rf._abc_6362_n4632), .Y(dp.rf._abc_6362_n3855) );
	NAND2X1 NAND2X1_3088 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4634) );
	NAND2X1 NAND2X1_3089 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<26>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4635) );
	NAND2X1 NAND2X1_3090 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4634), .B(dp.rf._abc_6362_n4635), .Y(dp.rf._abc_6362_n3856) );
	NAND2X1 NAND2X1_3091 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4637) );
	NAND2X1 NAND2X1_3092 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<27>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4638) );
	NAND2X1 NAND2X1_3093 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4637), .B(dp.rf._abc_6362_n4638), .Y(dp.rf._abc_6362_n3857) );
	NAND2X1 NAND2X1_3094 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4640) );
	NAND2X1 NAND2X1_3095 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<28>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4641) );
	NAND2X1 NAND2X1_3096 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4640), .B(dp.rf._abc_6362_n4641), .Y(dp.rf._abc_6362_n3858) );
	NAND2X1 NAND2X1_3097 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4643) );
	NAND2X1 NAND2X1_3098 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<29>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4644) );
	NAND2X1 NAND2X1_3099 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4643), .B(dp.rf._abc_6362_n4644), .Y(dp.rf._abc_6362_n3859) );
	NAND2X1 NAND2X1_3100 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4646) );
	NAND2X1 NAND2X1_3101 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<30>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4647) );
	NAND2X1 NAND2X1_3102 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4646), .B(dp.rf._abc_6362_n4647), .Y(dp.rf._abc_6362_n3860) );
	NAND2X1 NAND2X1_3103 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n4554), .Y(dp.rf._abc_6362_n4649) );
	NAND2X1 NAND2X1_3104 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_31_<31>), .B(dp.rf._abc_6362_n4556), .Y(dp.rf._abc_6362_n4650) );
	NAND2X1 NAND2X1_3105 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4649), .B(dp.rf._abc_6362_n4650), .Y(dp.rf._abc_6362_n3861) );
	NOR2X1 NOR2X1_217 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n3172_1), .Y(dp.rf._abc_6362_n4652) );
	NAND2X1 NAND2X1_3106 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4653) );
	INVX8 INVX8_30 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4654) );
	NAND2X1 NAND2X1_3107 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<0>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4655) );
	NAND2X1 NAND2X1_3108 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4653), .B(dp.rf._abc_6362_n4655), .Y(dp.rf._abc_6362_n3862) );
	NAND2X1 NAND2X1_3109 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4657) );
	NAND2X1 NAND2X1_3110 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<1>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4658) );
	NAND2X1 NAND2X1_3111 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4657), .B(dp.rf._abc_6362_n4658), .Y(dp.rf._abc_6362_n3863) );
	NAND2X1 NAND2X1_3112 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4660) );
	NAND2X1 NAND2X1_3113 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<2>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4661) );
	NAND2X1 NAND2X1_3114 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4660), .B(dp.rf._abc_6362_n4661), .Y(dp.rf._abc_6362_n3864) );
	NAND2X1 NAND2X1_3115 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4663) );
	NAND2X1 NAND2X1_3116 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<3>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4664) );
	NAND2X1 NAND2X1_3117 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4663), .B(dp.rf._abc_6362_n4664), .Y(dp.rf._abc_6362_n3865) );
	NAND2X1 NAND2X1_3118 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4666) );
	NAND2X1 NAND2X1_3119 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<4>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4667) );
	NAND2X1 NAND2X1_3120 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4666), .B(dp.rf._abc_6362_n4667), .Y(dp.rf._abc_6362_n3866) );
	NAND2X1 NAND2X1_3121 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4669) );
	NAND2X1 NAND2X1_3122 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<5>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4670) );
	NAND2X1 NAND2X1_3123 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4669), .B(dp.rf._abc_6362_n4670), .Y(dp.rf._abc_6362_n3867) );
	NAND2X1 NAND2X1_3124 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4672) );
	NAND2X1 NAND2X1_3125 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<6>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4673) );
	NAND2X1 NAND2X1_3126 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4672), .B(dp.rf._abc_6362_n4673), .Y(dp.rf._abc_6362_n3868) );
	NAND2X1 NAND2X1_3127 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4675) );
	NAND2X1 NAND2X1_3128 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<7>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4676) );
	NAND2X1 NAND2X1_3129 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4675), .B(dp.rf._abc_6362_n4676), .Y(dp.rf._abc_6362_n3869) );
	NAND2X1 NAND2X1_3130 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4678) );
	NAND2X1 NAND2X1_3131 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<8>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4679) );
	NAND2X1 NAND2X1_3132 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4678), .B(dp.rf._abc_6362_n4679), .Y(dp.rf._abc_6362_n3870) );
	NAND2X1 NAND2X1_3133 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4681) );
	NAND2X1 NAND2X1_3134 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<9>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4682) );
	NAND2X1 NAND2X1_3135 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4681), .B(dp.rf._abc_6362_n4682), .Y(dp.rf._abc_6362_n3871) );
	NAND2X1 NAND2X1_3136 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4684) );
	NAND2X1 NAND2X1_3137 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<10>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4685) );
	NAND2X1 NAND2X1_3138 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4684), .B(dp.rf._abc_6362_n4685), .Y(dp.rf._abc_6362_n3872) );
	NAND2X1 NAND2X1_3139 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4687) );
	NAND2X1 NAND2X1_3140 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<11>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4688) );
	NAND2X1 NAND2X1_3141 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4687), .B(dp.rf._abc_6362_n4688), .Y(dp.rf._abc_6362_n3873) );
	NAND2X1 NAND2X1_3142 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4690) );
	NAND2X1 NAND2X1_3143 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<12>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4691) );
	NAND2X1 NAND2X1_3144 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4690), .B(dp.rf._abc_6362_n4691), .Y(dp.rf._abc_6362_n3874) );
	NAND2X1 NAND2X1_3145 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4693) );
	NAND2X1 NAND2X1_3146 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<13>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4694) );
	NAND2X1 NAND2X1_3147 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4693), .B(dp.rf._abc_6362_n4694), .Y(dp.rf._abc_6362_n3875) );
	NAND2X1 NAND2X1_3148 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4696) );
	NAND2X1 NAND2X1_3149 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<14>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4697) );
	NAND2X1 NAND2X1_3150 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4696), .B(dp.rf._abc_6362_n4697), .Y(dp.rf._abc_6362_n3876) );
	NAND2X1 NAND2X1_3151 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4699) );
	NAND2X1 NAND2X1_3152 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<15>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4700) );
	NAND2X1 NAND2X1_3153 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4699), .B(dp.rf._abc_6362_n4700), .Y(dp.rf._abc_6362_n3877) );
	NAND2X1 NAND2X1_3154 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4702) );
	NAND2X1 NAND2X1_3155 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<16>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4703) );
	NAND2X1 NAND2X1_3156 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4702), .B(dp.rf._abc_6362_n4703), .Y(dp.rf._abc_6362_n3878) );
	NAND2X1 NAND2X1_3157 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4705) );
	NAND2X1 NAND2X1_3158 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<17>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4706) );
	NAND2X1 NAND2X1_3159 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4705), .B(dp.rf._abc_6362_n4706), .Y(dp.rf._abc_6362_n3879) );
	NAND2X1 NAND2X1_3160 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4708) );
	NAND2X1 NAND2X1_3161 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<18>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4709) );
	NAND2X1 NAND2X1_3162 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4708), .B(dp.rf._abc_6362_n4709), .Y(dp.rf._abc_6362_n3880) );
	NAND2X1 NAND2X1_3163 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4711) );
	NAND2X1 NAND2X1_3164 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<19>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4712) );
	NAND2X1 NAND2X1_3165 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4711), .B(dp.rf._abc_6362_n4712), .Y(dp.rf._abc_6362_n3881) );
	NAND2X1 NAND2X1_3166 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4714) );
	NAND2X1 NAND2X1_3167 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<20>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4715) );
	NAND2X1 NAND2X1_3168 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4714), .B(dp.rf._abc_6362_n4715), .Y(dp.rf._abc_6362_n3882) );
	NAND2X1 NAND2X1_3169 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4717) );
	NAND2X1 NAND2X1_3170 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<21>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4718) );
	NAND2X1 NAND2X1_3171 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4717), .B(dp.rf._abc_6362_n4718), .Y(dp.rf._abc_6362_n3883) );
	NAND2X1 NAND2X1_3172 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4720) );
	NAND2X1 NAND2X1_3173 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<22>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4721) );
	NAND2X1 NAND2X1_3174 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4720), .B(dp.rf._abc_6362_n4721), .Y(dp.rf._abc_6362_n3884) );
	NAND2X1 NAND2X1_3175 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4723) );
	NAND2X1 NAND2X1_3176 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<23>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4724) );
	NAND2X1 NAND2X1_3177 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4723), .B(dp.rf._abc_6362_n4724), .Y(dp.rf._abc_6362_n3885) );
	NAND2X1 NAND2X1_3178 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4726) );
	NAND2X1 NAND2X1_3179 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<24>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4727) );
	NAND2X1 NAND2X1_3180 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4726), .B(dp.rf._abc_6362_n4727), .Y(dp.rf._abc_6362_n3886) );
	NAND2X1 NAND2X1_3181 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4729) );
	NAND2X1 NAND2X1_3182 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<25>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4730) );
	NAND2X1 NAND2X1_3183 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4729), .B(dp.rf._abc_6362_n4730), .Y(dp.rf._abc_6362_n3887) );
	NAND2X1 NAND2X1_3184 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4732) );
	NAND2X1 NAND2X1_3185 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<26>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4733) );
	NAND2X1 NAND2X1_3186 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4732), .B(dp.rf._abc_6362_n4733), .Y(dp.rf._abc_6362_n3888) );
	NAND2X1 NAND2X1_3187 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4735) );
	NAND2X1 NAND2X1_3188 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<27>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4736) );
	NAND2X1 NAND2X1_3189 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4735), .B(dp.rf._abc_6362_n4736), .Y(dp.rf._abc_6362_n3889) );
	NAND2X1 NAND2X1_3190 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4738) );
	NAND2X1 NAND2X1_3191 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<28>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4739) );
	NAND2X1 NAND2X1_3192 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4738), .B(dp.rf._abc_6362_n4739), .Y(dp.rf._abc_6362_n3890) );
	NAND2X1 NAND2X1_3193 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4741) );
	NAND2X1 NAND2X1_3194 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<29>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4742) );
	NAND2X1 NAND2X1_3195 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4741), .B(dp.rf._abc_6362_n4742), .Y(dp.rf._abc_6362_n3891) );
	NAND2X1 NAND2X1_3196 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4744) );
	NAND2X1 NAND2X1_3197 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<30>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4745) );
	NAND2X1 NAND2X1_3198 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4744), .B(dp.rf._abc_6362_n4745), .Y(dp.rf._abc_6362_n3892) );
	NAND2X1 NAND2X1_3199 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n4652), .Y(dp.rf._abc_6362_n4747) );
	NAND2X1 NAND2X1_3200 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<31>), .B(dp.rf._abc_6362_n4654), .Y(dp.rf._abc_6362_n4748) );
	NAND2X1 NAND2X1_3201 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4747), .B(dp.rf._abc_6362_n4748), .Y(dp.rf._abc_6362_n3893) );
	NOR2X1 NOR2X1_218 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n3371_1), .Y(dp.rf._abc_6362_n4750) );
	NAND2X1 NAND2X1_3202 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4751) );
	INVX8 INVX8_31 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4752) );
	NAND2X1 NAND2X1_3203 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<0>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4753) );
	NAND2X1 NAND2X1_3204 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4751), .B(dp.rf._abc_6362_n4753), .Y(dp.rf._abc_6362_n3894) );
	NAND2X1 NAND2X1_3205 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4755) );
	NAND2X1 NAND2X1_3206 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<1>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4756) );
	NAND2X1 NAND2X1_3207 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4755), .B(dp.rf._abc_6362_n4756), .Y(dp.rf._abc_6362_n3895) );
	NAND2X1 NAND2X1_3208 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4758) );
	NAND2X1 NAND2X1_3209 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<2>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4759) );
	NAND2X1 NAND2X1_3210 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4758), .B(dp.rf._abc_6362_n4759), .Y(dp.rf._abc_6362_n3896) );
	NAND2X1 NAND2X1_3211 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4761) );
	NAND2X1 NAND2X1_3212 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<3>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4762) );
	NAND2X1 NAND2X1_3213 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4761), .B(dp.rf._abc_6362_n4762), .Y(dp.rf._abc_6362_n3897) );
	NAND2X1 NAND2X1_3214 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4764) );
	NAND2X1 NAND2X1_3215 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<4>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4765) );
	NAND2X1 NAND2X1_3216 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4764), .B(dp.rf._abc_6362_n4765), .Y(dp.rf._abc_6362_n3898) );
	NAND2X1 NAND2X1_3217 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4767) );
	NAND2X1 NAND2X1_3218 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<5>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4768) );
	NAND2X1 NAND2X1_3219 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4767), .B(dp.rf._abc_6362_n4768), .Y(dp.rf._abc_6362_n3899) );
	NAND2X1 NAND2X1_3220 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4770) );
	NAND2X1 NAND2X1_3221 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<6>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4771) );
	NAND2X1 NAND2X1_3222 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4770), .B(dp.rf._abc_6362_n4771), .Y(dp.rf._abc_6362_n3900) );
	NAND2X1 NAND2X1_3223 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4773) );
	NAND2X1 NAND2X1_3224 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<7>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4774) );
	NAND2X1 NAND2X1_3225 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4773), .B(dp.rf._abc_6362_n4774), .Y(dp.rf._abc_6362_n3901) );
	NAND2X1 NAND2X1_3226 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4776) );
	NAND2X1 NAND2X1_3227 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<8>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4777) );
	NAND2X1 NAND2X1_3228 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4776), .B(dp.rf._abc_6362_n4777), .Y(dp.rf._abc_6362_n3902) );
	NAND2X1 NAND2X1_3229 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4779) );
	NAND2X1 NAND2X1_3230 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<9>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4780) );
	NAND2X1 NAND2X1_3231 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4779), .B(dp.rf._abc_6362_n4780), .Y(dp.rf._abc_6362_n3903) );
	NAND2X1 NAND2X1_3232 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4782) );
	NAND2X1 NAND2X1_3233 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<10>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4783) );
	NAND2X1 NAND2X1_3234 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4782), .B(dp.rf._abc_6362_n4783), .Y(dp.rf._abc_6362_n3904) );
	NAND2X1 NAND2X1_3235 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4785) );
	NAND2X1 NAND2X1_3236 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<11>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4786) );
	NAND2X1 NAND2X1_3237 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4785), .B(dp.rf._abc_6362_n4786), .Y(dp.rf._abc_6362_n3905) );
	NAND2X1 NAND2X1_3238 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4788) );
	NAND2X1 NAND2X1_3239 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<12>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4789) );
	NAND2X1 NAND2X1_3240 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4788), .B(dp.rf._abc_6362_n4789), .Y(dp.rf._abc_6362_n3906) );
	NAND2X1 NAND2X1_3241 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4791) );
	NAND2X1 NAND2X1_3242 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<13>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4792) );
	NAND2X1 NAND2X1_3243 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4791), .B(dp.rf._abc_6362_n4792), .Y(dp.rf._abc_6362_n3907) );
	NAND2X1 NAND2X1_3244 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4794) );
	NAND2X1 NAND2X1_3245 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<14>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4795) );
	NAND2X1 NAND2X1_3246 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4794), .B(dp.rf._abc_6362_n4795), .Y(dp.rf._abc_6362_n3908) );
	NAND2X1 NAND2X1_3247 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4797) );
	NAND2X1 NAND2X1_3248 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<15>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4798) );
	NAND2X1 NAND2X1_3249 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4797), .B(dp.rf._abc_6362_n4798), .Y(dp.rf._abc_6362_n3909) );
	NAND2X1 NAND2X1_3250 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4800) );
	NAND2X1 NAND2X1_3251 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<16>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4801) );
	NAND2X1 NAND2X1_3252 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4800), .B(dp.rf._abc_6362_n4801), .Y(dp.rf._abc_6362_n3910) );
	NAND2X1 NAND2X1_3253 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4803) );
	NAND2X1 NAND2X1_3254 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<17>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4804) );
	NAND2X1 NAND2X1_3255 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4803), .B(dp.rf._abc_6362_n4804), .Y(dp.rf._abc_6362_n3911) );
	NAND2X1 NAND2X1_3256 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4806) );
	NAND2X1 NAND2X1_3257 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<18>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4807) );
	NAND2X1 NAND2X1_3258 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4806), .B(dp.rf._abc_6362_n4807), .Y(dp.rf._abc_6362_n3912) );
	NAND2X1 NAND2X1_3259 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4809) );
	NAND2X1 NAND2X1_3260 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<19>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4810) );
	NAND2X1 NAND2X1_3261 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4809), .B(dp.rf._abc_6362_n4810), .Y(dp.rf._abc_6362_n3913) );
	NAND2X1 NAND2X1_3262 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4812) );
	NAND2X1 NAND2X1_3263 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<20>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4813) );
	NAND2X1 NAND2X1_3264 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4812), .B(dp.rf._abc_6362_n4813), .Y(dp.rf._abc_6362_n3914) );
	NAND2X1 NAND2X1_3265 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4815) );
	NAND2X1 NAND2X1_3266 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<21>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4816) );
	NAND2X1 NAND2X1_3267 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4815), .B(dp.rf._abc_6362_n4816), .Y(dp.rf._abc_6362_n3915) );
	NAND2X1 NAND2X1_3268 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4818) );
	NAND2X1 NAND2X1_3269 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<22>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4819) );
	NAND2X1 NAND2X1_3270 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4818), .B(dp.rf._abc_6362_n4819), .Y(dp.rf._abc_6362_n3916) );
	NAND2X1 NAND2X1_3271 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4821) );
	NAND2X1 NAND2X1_3272 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<23>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4822) );
	NAND2X1 NAND2X1_3273 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4821), .B(dp.rf._abc_6362_n4822), .Y(dp.rf._abc_6362_n3917) );
	NAND2X1 NAND2X1_3274 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4824) );
	NAND2X1 NAND2X1_3275 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<24>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4825) );
	NAND2X1 NAND2X1_3276 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4824), .B(dp.rf._abc_6362_n4825), .Y(dp.rf._abc_6362_n3918) );
	NAND2X1 NAND2X1_3277 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4827) );
	NAND2X1 NAND2X1_3278 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<25>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4828) );
	NAND2X1 NAND2X1_3279 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4827), .B(dp.rf._abc_6362_n4828), .Y(dp.rf._abc_6362_n3919) );
	NAND2X1 NAND2X1_3280 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4830) );
	NAND2X1 NAND2X1_3281 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<26>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4831) );
	NAND2X1 NAND2X1_3282 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4830), .B(dp.rf._abc_6362_n4831), .Y(dp.rf._abc_6362_n3920) );
	NAND2X1 NAND2X1_3283 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4833) );
	NAND2X1 NAND2X1_3284 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<27>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4834) );
	NAND2X1 NAND2X1_3285 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4833), .B(dp.rf._abc_6362_n4834), .Y(dp.rf._abc_6362_n3921) );
	NAND2X1 NAND2X1_3286 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4836) );
	NAND2X1 NAND2X1_3287 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<28>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4837) );
	NAND2X1 NAND2X1_3288 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4836), .B(dp.rf._abc_6362_n4837), .Y(dp.rf._abc_6362_n3922) );
	NAND2X1 NAND2X1_3289 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4839) );
	NAND2X1 NAND2X1_3290 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<29>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4840) );
	NAND2X1 NAND2X1_3291 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4839), .B(dp.rf._abc_6362_n4840), .Y(dp.rf._abc_6362_n3923) );
	NAND2X1 NAND2X1_3292 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4842) );
	NAND2X1 NAND2X1_3293 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<30>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4843) );
	NAND2X1 NAND2X1_3294 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4842), .B(dp.rf._abc_6362_n4843), .Y(dp.rf._abc_6362_n3924) );
	NAND2X1 NAND2X1_3295 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n4750), .Y(dp.rf._abc_6362_n4845) );
	NAND2X1 NAND2X1_3296 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<31>), .B(dp.rf._abc_6362_n4752), .Y(dp.rf._abc_6362_n4846) );
	NAND2X1 NAND2X1_3297 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4845), .B(dp.rf._abc_6362_n4846), .Y(dp.rf._abc_6362_n3925) );
	NOR2X1 NOR2X1_219 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n3470_1), .Y(dp.rf._abc_6362_n4848) );
	NAND2X1 NAND2X1_3298 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4849) );
	INVX8 INVX8_32 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4850) );
	NAND2X1 NAND2X1_3299 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<0>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4851) );
	NAND2X1 NAND2X1_3300 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4849), .B(dp.rf._abc_6362_n4851), .Y(dp.rf._abc_6362_n3926) );
	NAND2X1 NAND2X1_3301 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4853) );
	NAND2X1 NAND2X1_3302 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<1>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4854) );
	NAND2X1 NAND2X1_3303 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4853), .B(dp.rf._abc_6362_n4854), .Y(dp.rf._abc_6362_n3927) );
	NAND2X1 NAND2X1_3304 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4856) );
	NAND2X1 NAND2X1_3305 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<2>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4857) );
	NAND2X1 NAND2X1_3306 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4856), .B(dp.rf._abc_6362_n4857), .Y(dp.rf._abc_6362_n3928) );
	NAND2X1 NAND2X1_3307 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4859) );
	NAND2X1 NAND2X1_3308 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<3>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4860) );
	NAND2X1 NAND2X1_3309 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4859), .B(dp.rf._abc_6362_n4860), .Y(dp.rf._abc_6362_n3929) );
	NAND2X1 NAND2X1_3310 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4862) );
	NAND2X1 NAND2X1_3311 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<4>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4863) );
	NAND2X1 NAND2X1_3312 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4862), .B(dp.rf._abc_6362_n4863), .Y(dp.rf._abc_6362_n3930) );
	NAND2X1 NAND2X1_3313 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4865) );
	NAND2X1 NAND2X1_3314 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<5>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4866) );
	NAND2X1 NAND2X1_3315 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4865), .B(dp.rf._abc_6362_n4866), .Y(dp.rf._abc_6362_n3931) );
	NAND2X1 NAND2X1_3316 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4868) );
	NAND2X1 NAND2X1_3317 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<6>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4869) );
	NAND2X1 NAND2X1_3318 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4868), .B(dp.rf._abc_6362_n4869), .Y(dp.rf._abc_6362_n3932) );
	NAND2X1 NAND2X1_3319 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4871) );
	NAND2X1 NAND2X1_3320 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<7>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4872) );
	NAND2X1 NAND2X1_3321 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4871), .B(dp.rf._abc_6362_n4872), .Y(dp.rf._abc_6362_n3933) );
	NAND2X1 NAND2X1_3322 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4874) );
	NAND2X1 NAND2X1_3323 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<8>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4875) );
	NAND2X1 NAND2X1_3324 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4874), .B(dp.rf._abc_6362_n4875), .Y(dp.rf._abc_6362_n3934) );
	NAND2X1 NAND2X1_3325 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4877) );
	NAND2X1 NAND2X1_3326 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<9>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4878) );
	NAND2X1 NAND2X1_3327 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4877), .B(dp.rf._abc_6362_n4878), .Y(dp.rf._abc_6362_n3935) );
	NAND2X1 NAND2X1_3328 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4880) );
	NAND2X1 NAND2X1_3329 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<10>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4881) );
	NAND2X1 NAND2X1_3330 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4880), .B(dp.rf._abc_6362_n4881), .Y(dp.rf._abc_6362_n3936) );
	NAND2X1 NAND2X1_3331 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4883) );
	NAND2X1 NAND2X1_3332 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<11>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4884) );
	NAND2X1 NAND2X1_3333 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4883), .B(dp.rf._abc_6362_n4884), .Y(dp.rf._abc_6362_n3937) );
	NAND2X1 NAND2X1_3334 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4886) );
	NAND2X1 NAND2X1_3335 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<12>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4887) );
	NAND2X1 NAND2X1_3336 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4886), .B(dp.rf._abc_6362_n4887), .Y(dp.rf._abc_6362_n3938) );
	NAND2X1 NAND2X1_3337 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4889) );
	NAND2X1 NAND2X1_3338 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<13>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4890) );
	NAND2X1 NAND2X1_3339 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4889), .B(dp.rf._abc_6362_n4890), .Y(dp.rf._abc_6362_n3939) );
	NAND2X1 NAND2X1_3340 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4892) );
	NAND2X1 NAND2X1_3341 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<14>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4893) );
	NAND2X1 NAND2X1_3342 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4892), .B(dp.rf._abc_6362_n4893), .Y(dp.rf._abc_6362_n3940) );
	NAND2X1 NAND2X1_3343 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4895) );
	NAND2X1 NAND2X1_3344 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<15>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4896) );
	NAND2X1 NAND2X1_3345 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4895), .B(dp.rf._abc_6362_n4896), .Y(dp.rf._abc_6362_n3941) );
	NAND2X1 NAND2X1_3346 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4898) );
	NAND2X1 NAND2X1_3347 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<16>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4899) );
	NAND2X1 NAND2X1_3348 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4898), .B(dp.rf._abc_6362_n4899), .Y(dp.rf._abc_6362_n3942) );
	NAND2X1 NAND2X1_3349 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4901) );
	NAND2X1 NAND2X1_3350 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<17>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4902) );
	NAND2X1 NAND2X1_3351 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4901), .B(dp.rf._abc_6362_n4902), .Y(dp.rf._abc_6362_n3943) );
	NAND2X1 NAND2X1_3352 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4904) );
	NAND2X1 NAND2X1_3353 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<18>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4905) );
	NAND2X1 NAND2X1_3354 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4904), .B(dp.rf._abc_6362_n4905), .Y(dp.rf._abc_6362_n3944) );
	NAND2X1 NAND2X1_3355 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4907) );
	NAND2X1 NAND2X1_3356 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<19>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4908) );
	NAND2X1 NAND2X1_3357 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4907), .B(dp.rf._abc_6362_n4908), .Y(dp.rf._abc_6362_n3945) );
	NAND2X1 NAND2X1_3358 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4910) );
	NAND2X1 NAND2X1_3359 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<20>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4911) );
	NAND2X1 NAND2X1_3360 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4910), .B(dp.rf._abc_6362_n4911), .Y(dp.rf._abc_6362_n3946) );
	NAND2X1 NAND2X1_3361 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4913) );
	NAND2X1 NAND2X1_3362 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<21>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4914) );
	NAND2X1 NAND2X1_3363 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4913), .B(dp.rf._abc_6362_n4914), .Y(dp.rf._abc_6362_n3947) );
	NAND2X1 NAND2X1_3364 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4916) );
	NAND2X1 NAND2X1_3365 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<22>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4917) );
	NAND2X1 NAND2X1_3366 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4916), .B(dp.rf._abc_6362_n4917), .Y(dp.rf._abc_6362_n3948) );
	NAND2X1 NAND2X1_3367 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4919) );
	NAND2X1 NAND2X1_3368 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<23>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4920) );
	NAND2X1 NAND2X1_3369 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4919), .B(dp.rf._abc_6362_n4920), .Y(dp.rf._abc_6362_n3949) );
	NAND2X1 NAND2X1_3370 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4922) );
	NAND2X1 NAND2X1_3371 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<24>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4923) );
	NAND2X1 NAND2X1_3372 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4922), .B(dp.rf._abc_6362_n4923), .Y(dp.rf._abc_6362_n3950) );
	NAND2X1 NAND2X1_3373 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4925) );
	NAND2X1 NAND2X1_3374 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<25>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4926) );
	NAND2X1 NAND2X1_3375 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4925), .B(dp.rf._abc_6362_n4926), .Y(dp.rf._abc_6362_n3951) );
	NAND2X1 NAND2X1_3376 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4928) );
	NAND2X1 NAND2X1_3377 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<26>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4929) );
	NAND2X1 NAND2X1_3378 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4928), .B(dp.rf._abc_6362_n4929), .Y(dp.rf._abc_6362_n3952) );
	NAND2X1 NAND2X1_3379 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4931) );
	NAND2X1 NAND2X1_3380 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<27>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4932) );
	NAND2X1 NAND2X1_3381 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4931), .B(dp.rf._abc_6362_n4932), .Y(dp.rf._abc_6362_n3953) );
	NAND2X1 NAND2X1_3382 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4934) );
	NAND2X1 NAND2X1_3383 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<28>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4935) );
	NAND2X1 NAND2X1_3384 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4934), .B(dp.rf._abc_6362_n4935), .Y(dp.rf._abc_6362_n3954) );
	NAND2X1 NAND2X1_3385 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4937) );
	NAND2X1 NAND2X1_3386 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<29>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4938) );
	NAND2X1 NAND2X1_3387 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4937), .B(dp.rf._abc_6362_n4938), .Y(dp.rf._abc_6362_n3955) );
	NAND2X1 NAND2X1_3388 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4940) );
	NAND2X1 NAND2X1_3389 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<30>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4941) );
	NAND2X1 NAND2X1_3390 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4940), .B(dp.rf._abc_6362_n4941), .Y(dp.rf._abc_6362_n3956) );
	NAND2X1 NAND2X1_3391 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n4848), .Y(dp.rf._abc_6362_n4943) );
	NAND2X1 NAND2X1_3392 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<31>), .B(dp.rf._abc_6362_n4850), .Y(dp.rf._abc_6362_n4944) );
	NAND2X1 NAND2X1_3393 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4943), .B(dp.rf._abc_6362_n4944), .Y(dp.rf._abc_6362_n3957) );
	NOR2X1 NOR2X1_220 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n3570_1), .Y(dp.rf._abc_6362_n4946) );
	NAND2X1 NAND2X1_3394 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4947) );
	INVX8 INVX8_33 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4948) );
	NAND2X1 NAND2X1_3395 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<0>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4949) );
	NAND2X1 NAND2X1_3396 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4947), .B(dp.rf._abc_6362_n4949), .Y(dp.rf._abc_6362_n3958) );
	NAND2X1 NAND2X1_3397 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4951) );
	NAND2X1 NAND2X1_3398 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<1>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4952) );
	NAND2X1 NAND2X1_3399 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4951), .B(dp.rf._abc_6362_n4952), .Y(dp.rf._abc_6362_n3959) );
	NAND2X1 NAND2X1_3400 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4954) );
	NAND2X1 NAND2X1_3401 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<2>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4955) );
	NAND2X1 NAND2X1_3402 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4954), .B(dp.rf._abc_6362_n4955), .Y(dp.rf._abc_6362_n3960) );
	NAND2X1 NAND2X1_3403 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4957) );
	NAND2X1 NAND2X1_3404 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<3>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4958) );
	NAND2X1 NAND2X1_3405 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4957), .B(dp.rf._abc_6362_n4958), .Y(dp.rf._abc_6362_n3961) );
	NAND2X1 NAND2X1_3406 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4960) );
	NAND2X1 NAND2X1_3407 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<4>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4961) );
	NAND2X1 NAND2X1_3408 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4960), .B(dp.rf._abc_6362_n4961), .Y(dp.rf._abc_6362_n3962) );
	NAND2X1 NAND2X1_3409 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4963) );
	NAND2X1 NAND2X1_3410 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<5>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4964) );
	NAND2X1 NAND2X1_3411 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4963), .B(dp.rf._abc_6362_n4964), .Y(dp.rf._abc_6362_n3963) );
	NAND2X1 NAND2X1_3412 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4966) );
	NAND2X1 NAND2X1_3413 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<6>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4967) );
	NAND2X1 NAND2X1_3414 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4966), .B(dp.rf._abc_6362_n4967), .Y(dp.rf._abc_6362_n3964) );
	NAND2X1 NAND2X1_3415 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4969) );
	NAND2X1 NAND2X1_3416 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<7>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4970) );
	NAND2X1 NAND2X1_3417 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4969), .B(dp.rf._abc_6362_n4970), .Y(dp.rf._abc_6362_n3965) );
	NAND2X1 NAND2X1_3418 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4972) );
	NAND2X1 NAND2X1_3419 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<8>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4973) );
	NAND2X1 NAND2X1_3420 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4972), .B(dp.rf._abc_6362_n4973), .Y(dp.rf._abc_6362_n3966) );
	NAND2X1 NAND2X1_3421 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4975) );
	NAND2X1 NAND2X1_3422 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<9>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4976) );
	NAND2X1 NAND2X1_3423 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4975), .B(dp.rf._abc_6362_n4976), .Y(dp.rf._abc_6362_n3967) );
	NAND2X1 NAND2X1_3424 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4978) );
	NAND2X1 NAND2X1_3425 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<10>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4979) );
	NAND2X1 NAND2X1_3426 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4978), .B(dp.rf._abc_6362_n4979), .Y(dp.rf._abc_6362_n3968) );
	NAND2X1 NAND2X1_3427 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4981) );
	NAND2X1 NAND2X1_3428 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<11>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4982) );
	NAND2X1 NAND2X1_3429 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4981), .B(dp.rf._abc_6362_n4982), .Y(dp.rf._abc_6362_n3969) );
	NAND2X1 NAND2X1_3430 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4984) );
	NAND2X1 NAND2X1_3431 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<12>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4985) );
	NAND2X1 NAND2X1_3432 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4984), .B(dp.rf._abc_6362_n4985), .Y(dp.rf._abc_6362_n3970) );
	NAND2X1 NAND2X1_3433 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4987) );
	NAND2X1 NAND2X1_3434 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<13>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4988) );
	NAND2X1 NAND2X1_3435 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4987), .B(dp.rf._abc_6362_n4988), .Y(dp.rf._abc_6362_n3971) );
	NAND2X1 NAND2X1_3436 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4990) );
	NAND2X1 NAND2X1_3437 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<14>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4991) );
	NAND2X1 NAND2X1_3438 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4990), .B(dp.rf._abc_6362_n4991), .Y(dp.rf._abc_6362_n3972) );
	NAND2X1 NAND2X1_3439 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4993) );
	NAND2X1 NAND2X1_3440 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<15>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4994) );
	NAND2X1 NAND2X1_3441 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4993), .B(dp.rf._abc_6362_n4994), .Y(dp.rf._abc_6362_n3973) );
	NAND2X1 NAND2X1_3442 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4996) );
	NAND2X1 NAND2X1_3443 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<16>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n4997) );
	NAND2X1 NAND2X1_3444 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4996), .B(dp.rf._abc_6362_n4997), .Y(dp.rf._abc_6362_n3974) );
	NAND2X1 NAND2X1_3445 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n4999) );
	NAND2X1 NAND2X1_3446 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<17>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5000) );
	NAND2X1 NAND2X1_3447 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n4999), .B(dp.rf._abc_6362_n5000), .Y(dp.rf._abc_6362_n3975) );
	NAND2X1 NAND2X1_3448 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5002) );
	NAND2X1 NAND2X1_3449 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<18>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5003) );
	NAND2X1 NAND2X1_3450 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5002), .B(dp.rf._abc_6362_n5003), .Y(dp.rf._abc_6362_n3976) );
	NAND2X1 NAND2X1_3451 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5005) );
	NAND2X1 NAND2X1_3452 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<19>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5006) );
	NAND2X1 NAND2X1_3453 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5005), .B(dp.rf._abc_6362_n5006), .Y(dp.rf._abc_6362_n3977) );
	NAND2X1 NAND2X1_3454 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5008) );
	NAND2X1 NAND2X1_3455 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<20>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5009) );
	NAND2X1 NAND2X1_3456 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5008), .B(dp.rf._abc_6362_n5009), .Y(dp.rf._abc_6362_n3978) );
	NAND2X1 NAND2X1_3457 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5011) );
	NAND2X1 NAND2X1_3458 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<21>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5012) );
	NAND2X1 NAND2X1_3459 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5011), .B(dp.rf._abc_6362_n5012), .Y(dp.rf._abc_6362_n3979) );
	NAND2X1 NAND2X1_3460 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5014) );
	NAND2X1 NAND2X1_3461 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<22>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5015) );
	NAND2X1 NAND2X1_3462 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5014), .B(dp.rf._abc_6362_n5015), .Y(dp.rf._abc_6362_n3980) );
	NAND2X1 NAND2X1_3463 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5017) );
	NAND2X1 NAND2X1_3464 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<23>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5018) );
	NAND2X1 NAND2X1_3465 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5017), .B(dp.rf._abc_6362_n5018), .Y(dp.rf._abc_6362_n3981) );
	NAND2X1 NAND2X1_3466 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5020) );
	NAND2X1 NAND2X1_3467 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<24>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5021) );
	NAND2X1 NAND2X1_3468 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5020), .B(dp.rf._abc_6362_n5021), .Y(dp.rf._abc_6362_n3982) );
	NAND2X1 NAND2X1_3469 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5023) );
	NAND2X1 NAND2X1_3470 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<25>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5024) );
	NAND2X1 NAND2X1_3471 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5023), .B(dp.rf._abc_6362_n5024), .Y(dp.rf._abc_6362_n3983) );
	NAND2X1 NAND2X1_3472 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5026) );
	NAND2X1 NAND2X1_3473 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<26>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5027) );
	NAND2X1 NAND2X1_3474 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5026), .B(dp.rf._abc_6362_n5027), .Y(dp.rf._abc_6362_n3984) );
	NAND2X1 NAND2X1_3475 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5029) );
	NAND2X1 NAND2X1_3476 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<27>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5030) );
	NAND2X1 NAND2X1_3477 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5029), .B(dp.rf._abc_6362_n5030), .Y(dp.rf._abc_6362_n3985) );
	NAND2X1 NAND2X1_3478 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5032) );
	NAND2X1 NAND2X1_3479 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<28>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5033) );
	NAND2X1 NAND2X1_3480 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5032), .B(dp.rf._abc_6362_n5033), .Y(dp.rf._abc_6362_n3986) );
	NAND2X1 NAND2X1_3481 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5035) );
	NAND2X1 NAND2X1_3482 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<29>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5036) );
	NAND2X1 NAND2X1_3483 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5035), .B(dp.rf._abc_6362_n5036), .Y(dp.rf._abc_6362_n3987) );
	NAND2X1 NAND2X1_3484 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5038) );
	NAND2X1 NAND2X1_3485 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<30>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5039) );
	NAND2X1 NAND2X1_3486 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5038), .B(dp.rf._abc_6362_n5039), .Y(dp.rf._abc_6362_n3988) );
	NAND2X1 NAND2X1_3487 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n4946), .Y(dp.rf._abc_6362_n5041) );
	NAND2X1 NAND2X1_3488 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<31>), .B(dp.rf._abc_6362_n4948), .Y(dp.rf._abc_6362_n5042) );
	NAND2X1 NAND2X1_3489 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5041), .B(dp.rf._abc_6362_n5042), .Y(dp.rf._abc_6362_n3989) );
	NOR2X1 NOR2X1_221 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n3669_1), .Y(dp.rf._abc_6362_n5044) );
	NAND2X1 NAND2X1_3490 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5045) );
	INVX8 INVX8_34 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5046) );
	NAND2X1 NAND2X1_3491 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<0>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5047) );
	NAND2X1 NAND2X1_3492 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5045), .B(dp.rf._abc_6362_n5047), .Y(dp.rf._abc_6362_n3990) );
	NAND2X1 NAND2X1_3493 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5049) );
	NAND2X1 NAND2X1_3494 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<1>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5050) );
	NAND2X1 NAND2X1_3495 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5049), .B(dp.rf._abc_6362_n5050), .Y(dp.rf._abc_6362_n3991) );
	NAND2X1 NAND2X1_3496 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5052) );
	NAND2X1 NAND2X1_3497 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<2>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5053) );
	NAND2X1 NAND2X1_3498 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5052), .B(dp.rf._abc_6362_n5053), .Y(dp.rf._abc_6362_n3992) );
	NAND2X1 NAND2X1_3499 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5055) );
	NAND2X1 NAND2X1_3500 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<3>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5056) );
	NAND2X1 NAND2X1_3501 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5055), .B(dp.rf._abc_6362_n5056), .Y(dp.rf._abc_6362_n3993) );
	NAND2X1 NAND2X1_3502 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5058) );
	NAND2X1 NAND2X1_3503 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<4>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5059) );
	NAND2X1 NAND2X1_3504 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5058), .B(dp.rf._abc_6362_n5059), .Y(dp.rf._abc_6362_n3994) );
	NAND2X1 NAND2X1_3505 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5061) );
	NAND2X1 NAND2X1_3506 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<5>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5062) );
	NAND2X1 NAND2X1_3507 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5061), .B(dp.rf._abc_6362_n5062), .Y(dp.rf._abc_6362_n3995) );
	NAND2X1 NAND2X1_3508 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5064) );
	NAND2X1 NAND2X1_3509 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<6>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5065) );
	NAND2X1 NAND2X1_3510 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5064), .B(dp.rf._abc_6362_n5065), .Y(dp.rf._abc_6362_n3996) );
	NAND2X1 NAND2X1_3511 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5067) );
	NAND2X1 NAND2X1_3512 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<7>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5068) );
	NAND2X1 NAND2X1_3513 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5067), .B(dp.rf._abc_6362_n5068), .Y(dp.rf._abc_6362_n3997) );
	NAND2X1 NAND2X1_3514 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5070) );
	NAND2X1 NAND2X1_3515 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<8>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5071) );
	NAND2X1 NAND2X1_3516 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5070), .B(dp.rf._abc_6362_n5071), .Y(dp.rf._abc_6362_n3998) );
	NAND2X1 NAND2X1_3517 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5073) );
	NAND2X1 NAND2X1_3518 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<9>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5074) );
	NAND2X1 NAND2X1_3519 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5073), .B(dp.rf._abc_6362_n5074), .Y(dp.rf._abc_6362_n3999) );
	NAND2X1 NAND2X1_3520 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5076) );
	NAND2X1 NAND2X1_3521 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<10>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5077) );
	NAND2X1 NAND2X1_3522 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5076), .B(dp.rf._abc_6362_n5077), .Y(dp.rf._abc_6362_n4000) );
	NAND2X1 NAND2X1_3523 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5079) );
	NAND2X1 NAND2X1_3524 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<11>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5080) );
	NAND2X1 NAND2X1_3525 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5079), .B(dp.rf._abc_6362_n5080), .Y(dp.rf._abc_6362_n4001) );
	NAND2X1 NAND2X1_3526 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5082) );
	NAND2X1 NAND2X1_3527 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<12>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5083) );
	NAND2X1 NAND2X1_3528 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5082), .B(dp.rf._abc_6362_n5083), .Y(dp.rf._abc_6362_n4002) );
	NAND2X1 NAND2X1_3529 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5085) );
	NAND2X1 NAND2X1_3530 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<13>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5086) );
	NAND2X1 NAND2X1_3531 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5085), .B(dp.rf._abc_6362_n5086), .Y(dp.rf._abc_6362_n4003) );
	NAND2X1 NAND2X1_3532 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5088) );
	NAND2X1 NAND2X1_3533 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<14>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5089) );
	NAND2X1 NAND2X1_3534 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5088), .B(dp.rf._abc_6362_n5089), .Y(dp.rf._abc_6362_n4004) );
	NAND2X1 NAND2X1_3535 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5091) );
	NAND2X1 NAND2X1_3536 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<15>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5092) );
	NAND2X1 NAND2X1_3537 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5091), .B(dp.rf._abc_6362_n5092), .Y(dp.rf._abc_6362_n4005) );
	NAND2X1 NAND2X1_3538 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5094) );
	NAND2X1 NAND2X1_3539 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<16>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5095) );
	NAND2X1 NAND2X1_3540 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5094), .B(dp.rf._abc_6362_n5095), .Y(dp.rf._abc_6362_n4006) );
	NAND2X1 NAND2X1_3541 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5097) );
	NAND2X1 NAND2X1_3542 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<17>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5098) );
	NAND2X1 NAND2X1_3543 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5097), .B(dp.rf._abc_6362_n5098), .Y(dp.rf._abc_6362_n4007) );
	NAND2X1 NAND2X1_3544 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5100) );
	NAND2X1 NAND2X1_3545 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<18>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5101) );
	NAND2X1 NAND2X1_3546 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5100), .B(dp.rf._abc_6362_n5101), .Y(dp.rf._abc_6362_n4008) );
	NAND2X1 NAND2X1_3547 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5103) );
	NAND2X1 NAND2X1_3548 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<19>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5104) );
	NAND2X1 NAND2X1_3549 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5103), .B(dp.rf._abc_6362_n5104), .Y(dp.rf._abc_6362_n4009) );
	NAND2X1 NAND2X1_3550 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5106) );
	NAND2X1 NAND2X1_3551 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<20>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5107) );
	NAND2X1 NAND2X1_3552 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5106), .B(dp.rf._abc_6362_n5107), .Y(dp.rf._abc_6362_n4010) );
	NAND2X1 NAND2X1_3553 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5109) );
	NAND2X1 NAND2X1_3554 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<21>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5110) );
	NAND2X1 NAND2X1_3555 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5109), .B(dp.rf._abc_6362_n5110), .Y(dp.rf._abc_6362_n4011) );
	NAND2X1 NAND2X1_3556 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5112) );
	NAND2X1 NAND2X1_3557 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<22>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5113) );
	NAND2X1 NAND2X1_3558 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5112), .B(dp.rf._abc_6362_n5113), .Y(dp.rf._abc_6362_n4012) );
	NAND2X1 NAND2X1_3559 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5115) );
	NAND2X1 NAND2X1_3560 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<23>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5116) );
	NAND2X1 NAND2X1_3561 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5115), .B(dp.rf._abc_6362_n5116), .Y(dp.rf._abc_6362_n4013) );
	NAND2X1 NAND2X1_3562 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5118) );
	NAND2X1 NAND2X1_3563 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<24>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5119) );
	NAND2X1 NAND2X1_3564 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5118), .B(dp.rf._abc_6362_n5119), .Y(dp.rf._abc_6362_n4014) );
	NAND2X1 NAND2X1_3565 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5121) );
	NAND2X1 NAND2X1_3566 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<25>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5122) );
	NAND2X1 NAND2X1_3567 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5121), .B(dp.rf._abc_6362_n5122), .Y(dp.rf._abc_6362_n4015) );
	NAND2X1 NAND2X1_3568 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5124) );
	NAND2X1 NAND2X1_3569 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<26>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5125) );
	NAND2X1 NAND2X1_3570 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5124), .B(dp.rf._abc_6362_n5125), .Y(dp.rf._abc_6362_n4016) );
	NAND2X1 NAND2X1_3571 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5127) );
	NAND2X1 NAND2X1_3572 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<27>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5128) );
	NAND2X1 NAND2X1_3573 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5127), .B(dp.rf._abc_6362_n5128), .Y(dp.rf._abc_6362_n4017) );
	NAND2X1 NAND2X1_3574 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5130) );
	NAND2X1 NAND2X1_3575 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<28>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5131) );
	NAND2X1 NAND2X1_3576 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5130), .B(dp.rf._abc_6362_n5131), .Y(dp.rf._abc_6362_n4018) );
	NAND2X1 NAND2X1_3577 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5133) );
	NAND2X1 NAND2X1_3578 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<29>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5134) );
	NAND2X1 NAND2X1_3579 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5133), .B(dp.rf._abc_6362_n5134), .Y(dp.rf._abc_6362_n4019) );
	NAND2X1 NAND2X1_3580 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5136) );
	NAND2X1 NAND2X1_3581 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<30>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5137) );
	NAND2X1 NAND2X1_3582 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5136), .B(dp.rf._abc_6362_n5137), .Y(dp.rf._abc_6362_n4020) );
	NAND2X1 NAND2X1_3583 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n5044), .Y(dp.rf._abc_6362_n5139) );
	NAND2X1 NAND2X1_3584 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<31>), .B(dp.rf._abc_6362_n5046), .Y(dp.rf._abc_6362_n5140) );
	NAND2X1 NAND2X1_3585 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5139), .B(dp.rf._abc_6362_n5140), .Y(dp.rf._abc_6362_n4021) );
	NOR2X1 NOR2X1_222 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n3768_1), .Y(dp.rf._abc_6362_n5142) );
	NAND2X1 NAND2X1_3586 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5143) );
	INVX8 INVX8_35 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5144) );
	NAND2X1 NAND2X1_3587 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<0>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5145) );
	NAND2X1 NAND2X1_3588 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5143), .B(dp.rf._abc_6362_n5145), .Y(dp.rf._abc_6362_n4022) );
	NAND2X1 NAND2X1_3589 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5147) );
	NAND2X1 NAND2X1_3590 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<1>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5148) );
	NAND2X1 NAND2X1_3591 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5147), .B(dp.rf._abc_6362_n5148), .Y(dp.rf._abc_6362_n4023) );
	NAND2X1 NAND2X1_3592 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5150) );
	NAND2X1 NAND2X1_3593 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<2>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5151) );
	NAND2X1 NAND2X1_3594 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5150), .B(dp.rf._abc_6362_n5151), .Y(dp.rf._abc_6362_n4024) );
	NAND2X1 NAND2X1_3595 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5153) );
	NAND2X1 NAND2X1_3596 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<3>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5154) );
	NAND2X1 NAND2X1_3597 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5153), .B(dp.rf._abc_6362_n5154), .Y(dp.rf._abc_6362_n4025) );
	NAND2X1 NAND2X1_3598 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5156) );
	NAND2X1 NAND2X1_3599 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<4>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5157) );
	NAND2X1 NAND2X1_3600 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5156), .B(dp.rf._abc_6362_n5157), .Y(dp.rf._abc_6362_n4026) );
	NAND2X1 NAND2X1_3601 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5159) );
	NAND2X1 NAND2X1_3602 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<5>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5160) );
	NAND2X1 NAND2X1_3603 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5159), .B(dp.rf._abc_6362_n5160), .Y(dp.rf._abc_6362_n4027) );
	NAND2X1 NAND2X1_3604 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5162) );
	NAND2X1 NAND2X1_3605 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<6>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5163) );
	NAND2X1 NAND2X1_3606 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5162), .B(dp.rf._abc_6362_n5163), .Y(dp.rf._abc_6362_n4028) );
	NAND2X1 NAND2X1_3607 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5165) );
	NAND2X1 NAND2X1_3608 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<7>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5166) );
	NAND2X1 NAND2X1_3609 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5165), .B(dp.rf._abc_6362_n5166), .Y(dp.rf._abc_6362_n4029) );
	NAND2X1 NAND2X1_3610 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5168) );
	NAND2X1 NAND2X1_3611 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<8>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5169) );
	NAND2X1 NAND2X1_3612 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5168), .B(dp.rf._abc_6362_n5169), .Y(dp.rf._abc_6362_n4030) );
	NAND2X1 NAND2X1_3613 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5171) );
	NAND2X1 NAND2X1_3614 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<9>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5172) );
	NAND2X1 NAND2X1_3615 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5171), .B(dp.rf._abc_6362_n5172), .Y(dp.rf._abc_6362_n4031) );
	NAND2X1 NAND2X1_3616 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5174) );
	NAND2X1 NAND2X1_3617 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<10>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5175) );
	NAND2X1 NAND2X1_3618 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5174), .B(dp.rf._abc_6362_n5175), .Y(dp.rf._abc_6362_n4032) );
	NAND2X1 NAND2X1_3619 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5177) );
	NAND2X1 NAND2X1_3620 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<11>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5178) );
	NAND2X1 NAND2X1_3621 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5177), .B(dp.rf._abc_6362_n5178), .Y(dp.rf._abc_6362_n4033) );
	NAND2X1 NAND2X1_3622 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5180) );
	NAND2X1 NAND2X1_3623 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<12>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5181) );
	NAND2X1 NAND2X1_3624 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5180), .B(dp.rf._abc_6362_n5181), .Y(dp.rf._abc_6362_n4034) );
	NAND2X1 NAND2X1_3625 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5183) );
	NAND2X1 NAND2X1_3626 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<13>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5184) );
	NAND2X1 NAND2X1_3627 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5183), .B(dp.rf._abc_6362_n5184), .Y(dp.rf._abc_6362_n4035) );
	NAND2X1 NAND2X1_3628 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5186) );
	NAND2X1 NAND2X1_3629 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<14>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5187) );
	NAND2X1 NAND2X1_3630 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5186), .B(dp.rf._abc_6362_n5187), .Y(dp.rf._abc_6362_n4036) );
	NAND2X1 NAND2X1_3631 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5189) );
	NAND2X1 NAND2X1_3632 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<15>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5190) );
	NAND2X1 NAND2X1_3633 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5189), .B(dp.rf._abc_6362_n5190), .Y(dp.rf._abc_6362_n4037) );
	NAND2X1 NAND2X1_3634 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5192) );
	NAND2X1 NAND2X1_3635 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<16>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5193) );
	NAND2X1 NAND2X1_3636 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5192), .B(dp.rf._abc_6362_n5193), .Y(dp.rf._abc_6362_n4038) );
	NAND2X1 NAND2X1_3637 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5195) );
	NAND2X1 NAND2X1_3638 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<17>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5196) );
	NAND2X1 NAND2X1_3639 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5195), .B(dp.rf._abc_6362_n5196), .Y(dp.rf._abc_6362_n4039) );
	NAND2X1 NAND2X1_3640 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5198) );
	NAND2X1 NAND2X1_3641 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<18>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5199) );
	NAND2X1 NAND2X1_3642 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5198), .B(dp.rf._abc_6362_n5199), .Y(dp.rf._abc_6362_n4040) );
	NAND2X1 NAND2X1_3643 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5201) );
	NAND2X1 NAND2X1_3644 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<19>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5202) );
	NAND2X1 NAND2X1_3645 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5201), .B(dp.rf._abc_6362_n5202), .Y(dp.rf._abc_6362_n4041) );
	NAND2X1 NAND2X1_3646 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5204) );
	NAND2X1 NAND2X1_3647 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<20>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5205) );
	NAND2X1 NAND2X1_3648 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5204), .B(dp.rf._abc_6362_n5205), .Y(dp.rf._abc_6362_n4042) );
	NAND2X1 NAND2X1_3649 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5207) );
	NAND2X1 NAND2X1_3650 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<21>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5208) );
	NAND2X1 NAND2X1_3651 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5207), .B(dp.rf._abc_6362_n5208), .Y(dp.rf._abc_6362_n4043) );
	NAND2X1 NAND2X1_3652 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5210) );
	NAND2X1 NAND2X1_3653 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<22>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5211) );
	NAND2X1 NAND2X1_3654 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5210), .B(dp.rf._abc_6362_n5211), .Y(dp.rf._abc_6362_n4044) );
	NAND2X1 NAND2X1_3655 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5213) );
	NAND2X1 NAND2X1_3656 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<23>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5214) );
	NAND2X1 NAND2X1_3657 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5213), .B(dp.rf._abc_6362_n5214), .Y(dp.rf._abc_6362_n4045) );
	NAND2X1 NAND2X1_3658 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5216) );
	NAND2X1 NAND2X1_3659 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<24>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5217) );
	NAND2X1 NAND2X1_3660 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5216), .B(dp.rf._abc_6362_n5217), .Y(dp.rf._abc_6362_n4046) );
	NAND2X1 NAND2X1_3661 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5219) );
	NAND2X1 NAND2X1_3662 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<25>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5220) );
	NAND2X1 NAND2X1_3663 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5219), .B(dp.rf._abc_6362_n5220), .Y(dp.rf._abc_6362_n4047) );
	NAND2X1 NAND2X1_3664 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5222) );
	NAND2X1 NAND2X1_3665 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<26>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5223) );
	NAND2X1 NAND2X1_3666 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5222), .B(dp.rf._abc_6362_n5223), .Y(dp.rf._abc_6362_n4048) );
	NAND2X1 NAND2X1_3667 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5225) );
	NAND2X1 NAND2X1_3668 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<27>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5226) );
	NAND2X1 NAND2X1_3669 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5225), .B(dp.rf._abc_6362_n5226), .Y(dp.rf._abc_6362_n4049) );
	NAND2X1 NAND2X1_3670 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5228) );
	NAND2X1 NAND2X1_3671 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<28>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5229) );
	NAND2X1 NAND2X1_3672 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5228), .B(dp.rf._abc_6362_n5229), .Y(dp.rf._abc_6362_n4050) );
	NAND2X1 NAND2X1_3673 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5231) );
	NAND2X1 NAND2X1_3674 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<29>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5232) );
	NAND2X1 NAND2X1_3675 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5231), .B(dp.rf._abc_6362_n5232), .Y(dp.rf._abc_6362_n4051) );
	NAND2X1 NAND2X1_3676 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5234) );
	NAND2X1 NAND2X1_3677 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<30>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5235) );
	NAND2X1 NAND2X1_3678 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5234), .B(dp.rf._abc_6362_n5235), .Y(dp.rf._abc_6362_n4052) );
	NAND2X1 NAND2X1_3679 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n5142), .Y(dp.rf._abc_6362_n5237) );
	NAND2X1 NAND2X1_3680 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<31>), .B(dp.rf._abc_6362_n5144), .Y(dp.rf._abc_6362_n5238) );
	NAND2X1 NAND2X1_3681 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5237), .B(dp.rf._abc_6362_n5238), .Y(dp.rf._abc_6362_n4053) );
	NOR2X1 NOR2X1_223 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n2162), .B(dp.rf._abc_6362_n3867_1), .Y(dp.rf._abc_6362_n5240) );
	NAND2X1 NAND2X1_3682 ( .gnd(gnd), .vdd(vdd), .A(dp.result_0_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5241) );
	INVX8 INVX8_36 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5242) );
	NAND2X1 NAND2X1_3683 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<0>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5243) );
	NAND2X1 NAND2X1_3684 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5241), .B(dp.rf._abc_6362_n5243), .Y(dp.rf._abc_6362_n4054) );
	NAND2X1 NAND2X1_3685 ( .gnd(gnd), .vdd(vdd), .A(dp.result_1_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5245) );
	NAND2X1 NAND2X1_3686 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<1>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5246) );
	NAND2X1 NAND2X1_3687 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5245), .B(dp.rf._abc_6362_n5246), .Y(dp.rf._abc_6362_n4055) );
	NAND2X1 NAND2X1_3688 ( .gnd(gnd), .vdd(vdd), .A(dp.result_2_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5248) );
	NAND2X1 NAND2X1_3689 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<2>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5249) );
	NAND2X1 NAND2X1_3690 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5248), .B(dp.rf._abc_6362_n5249), .Y(dp.rf._abc_6362_n4056) );
	NAND2X1 NAND2X1_3691 ( .gnd(gnd), .vdd(vdd), .A(dp.result_3_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5251) );
	NAND2X1 NAND2X1_3692 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<3>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5252) );
	NAND2X1 NAND2X1_3693 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5251), .B(dp.rf._abc_6362_n5252), .Y(dp.rf._abc_6362_n4057) );
	NAND2X1 NAND2X1_3694 ( .gnd(gnd), .vdd(vdd), .A(dp.result_4_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5254) );
	NAND2X1 NAND2X1_3695 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<4>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5255) );
	NAND2X1 NAND2X1_3696 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5254), .B(dp.rf._abc_6362_n5255), .Y(dp.rf._abc_6362_n4058) );
	NAND2X1 NAND2X1_3697 ( .gnd(gnd), .vdd(vdd), .A(dp.result_5_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5257) );
	NAND2X1 NAND2X1_3698 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<5>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5258) );
	NAND2X1 NAND2X1_3699 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5257), .B(dp.rf._abc_6362_n5258), .Y(dp.rf._abc_6362_n4059) );
	NAND2X1 NAND2X1_3700 ( .gnd(gnd), .vdd(vdd), .A(dp.result_6_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5260) );
	NAND2X1 NAND2X1_3701 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<6>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5261) );
	NAND2X1 NAND2X1_3702 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5260), .B(dp.rf._abc_6362_n5261), .Y(dp.rf._abc_6362_n4060) );
	NAND2X1 NAND2X1_3703 ( .gnd(gnd), .vdd(vdd), .A(dp.result_7_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5263) );
	NAND2X1 NAND2X1_3704 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<7>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5264) );
	NAND2X1 NAND2X1_3705 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5263), .B(dp.rf._abc_6362_n5264), .Y(dp.rf._abc_6362_n4061) );
	NAND2X1 NAND2X1_3706 ( .gnd(gnd), .vdd(vdd), .A(dp.result_8_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5266) );
	NAND2X1 NAND2X1_3707 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<8>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5267) );
	NAND2X1 NAND2X1_3708 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5266), .B(dp.rf._abc_6362_n5267), .Y(dp.rf._abc_6362_n4062) );
	NAND2X1 NAND2X1_3709 ( .gnd(gnd), .vdd(vdd), .A(dp.result_9_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5269) );
	NAND2X1 NAND2X1_3710 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<9>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5270) );
	NAND2X1 NAND2X1_3711 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5269), .B(dp.rf._abc_6362_n5270), .Y(dp.rf._abc_6362_n4063) );
	NAND2X1 NAND2X1_3712 ( .gnd(gnd), .vdd(vdd), .A(dp.result_10_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5272) );
	NAND2X1 NAND2X1_3713 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<10>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5273) );
	NAND2X1 NAND2X1_3714 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5272), .B(dp.rf._abc_6362_n5273), .Y(dp.rf._abc_6362_n4064) );
	NAND2X1 NAND2X1_3715 ( .gnd(gnd), .vdd(vdd), .A(dp.result_11_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5275) );
	NAND2X1 NAND2X1_3716 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<11>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5276) );
	NAND2X1 NAND2X1_3717 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5275), .B(dp.rf._abc_6362_n5276), .Y(dp.rf._abc_6362_n4065) );
	NAND2X1 NAND2X1_3718 ( .gnd(gnd), .vdd(vdd), .A(dp.result_12_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5278) );
	NAND2X1 NAND2X1_3719 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<12>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5279) );
	NAND2X1 NAND2X1_3720 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5278), .B(dp.rf._abc_6362_n5279), .Y(dp.rf._abc_6362_n4066) );
	NAND2X1 NAND2X1_3721 ( .gnd(gnd), .vdd(vdd), .A(dp.result_13_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5281) );
	NAND2X1 NAND2X1_3722 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<13>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5282) );
	NAND2X1 NAND2X1_3723 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5281), .B(dp.rf._abc_6362_n5282), .Y(dp.rf._abc_6362_n4067) );
	NAND2X1 NAND2X1_3724 ( .gnd(gnd), .vdd(vdd), .A(dp.result_14_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5284) );
	NAND2X1 NAND2X1_3725 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<14>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5285) );
	NAND2X1 NAND2X1_3726 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5284), .B(dp.rf._abc_6362_n5285), .Y(dp.rf._abc_6362_n4068) );
	NAND2X1 NAND2X1_3727 ( .gnd(gnd), .vdd(vdd), .A(dp.result_15_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5287) );
	NAND2X1 NAND2X1_3728 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<15>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5288) );
	NAND2X1 NAND2X1_3729 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5287), .B(dp.rf._abc_6362_n5288), .Y(dp.rf._abc_6362_n4069) );
	NAND2X1 NAND2X1_3730 ( .gnd(gnd), .vdd(vdd), .A(dp.result_16_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5290) );
	NAND2X1 NAND2X1_3731 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<16>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5291) );
	NAND2X1 NAND2X1_3732 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5290), .B(dp.rf._abc_6362_n5291), .Y(dp.rf._abc_6362_n4070) );
	NAND2X1 NAND2X1_3733 ( .gnd(gnd), .vdd(vdd), .A(dp.result_17_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5293) );
	NAND2X1 NAND2X1_3734 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<17>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5294) );
	NAND2X1 NAND2X1_3735 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5293), .B(dp.rf._abc_6362_n5294), .Y(dp.rf._abc_6362_n4071) );
	NAND2X1 NAND2X1_3736 ( .gnd(gnd), .vdd(vdd), .A(dp.result_18_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5296) );
	NAND2X1 NAND2X1_3737 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<18>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5297) );
	NAND2X1 NAND2X1_3738 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5296), .B(dp.rf._abc_6362_n5297), .Y(dp.rf._abc_6362_n4072) );
	NAND2X1 NAND2X1_3739 ( .gnd(gnd), .vdd(vdd), .A(dp.result_19_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5299) );
	NAND2X1 NAND2X1_3740 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<19>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5300) );
	NAND2X1 NAND2X1_3741 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5299), .B(dp.rf._abc_6362_n5300), .Y(dp.rf._abc_6362_n4073) );
	NAND2X1 NAND2X1_3742 ( .gnd(gnd), .vdd(vdd), .A(dp.result_20_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5302) );
	NAND2X1 NAND2X1_3743 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<20>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5303) );
	NAND2X1 NAND2X1_3744 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5302), .B(dp.rf._abc_6362_n5303), .Y(dp.rf._abc_6362_n4074) );
	NAND2X1 NAND2X1_3745 ( .gnd(gnd), .vdd(vdd), .A(dp.result_21_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5305) );
	NAND2X1 NAND2X1_3746 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<21>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5306) );
	NAND2X1 NAND2X1_3747 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5305), .B(dp.rf._abc_6362_n5306), .Y(dp.rf._abc_6362_n4075) );
	NAND2X1 NAND2X1_3748 ( .gnd(gnd), .vdd(vdd), .A(dp.result_22_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5308) );
	NAND2X1 NAND2X1_3749 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<22>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5309) );
	NAND2X1 NAND2X1_3750 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5308), .B(dp.rf._abc_6362_n5309), .Y(dp.rf._abc_6362_n4076) );
	NAND2X1 NAND2X1_3751 ( .gnd(gnd), .vdd(vdd), .A(dp.result_23_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5311) );
	NAND2X1 NAND2X1_3752 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<23>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5312) );
	NAND2X1 NAND2X1_3753 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5311), .B(dp.rf._abc_6362_n5312), .Y(dp.rf._abc_6362_n4077) );
	NAND2X1 NAND2X1_3754 ( .gnd(gnd), .vdd(vdd), .A(dp.result_24_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5314) );
	NAND2X1 NAND2X1_3755 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<24>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5315) );
	NAND2X1 NAND2X1_3756 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5314), .B(dp.rf._abc_6362_n5315), .Y(dp.rf._abc_6362_n4078) );
	NAND2X1 NAND2X1_3757 ( .gnd(gnd), .vdd(vdd), .A(dp.result_25_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5317) );
	NAND2X1 NAND2X1_3758 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<25>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5318) );
	NAND2X1 NAND2X1_3759 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5317), .B(dp.rf._abc_6362_n5318), .Y(dp.rf._abc_6362_n4079) );
	NAND2X1 NAND2X1_3760 ( .gnd(gnd), .vdd(vdd), .A(dp.result_26_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5320) );
	NAND2X1 NAND2X1_3761 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<26>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5321) );
	NAND2X1 NAND2X1_3762 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5320), .B(dp.rf._abc_6362_n5321), .Y(dp.rf._abc_6362_n4080) );
	NAND2X1 NAND2X1_3763 ( .gnd(gnd), .vdd(vdd), .A(dp.result_27_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5323) );
	NAND2X1 NAND2X1_3764 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<27>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5324) );
	NAND2X1 NAND2X1_3765 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5323), .B(dp.rf._abc_6362_n5324), .Y(dp.rf._abc_6362_n4081) );
	NAND2X1 NAND2X1_3766 ( .gnd(gnd), .vdd(vdd), .A(dp.result_28_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5326) );
	NAND2X1 NAND2X1_3767 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<28>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5327) );
	NAND2X1 NAND2X1_3768 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5326), .B(dp.rf._abc_6362_n5327), .Y(dp.rf._abc_6362_n4082) );
	NAND2X1 NAND2X1_3769 ( .gnd(gnd), .vdd(vdd), .A(dp.result_29_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5329) );
	NAND2X1 NAND2X1_3770 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<29>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5330) );
	NAND2X1 NAND2X1_3771 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5329), .B(dp.rf._abc_6362_n5330), .Y(dp.rf._abc_6362_n4083) );
	NAND2X1 NAND2X1_3772 ( .gnd(gnd), .vdd(vdd), .A(dp.result_30_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5332) );
	NAND2X1 NAND2X1_3773 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<30>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5333) );
	NAND2X1 NAND2X1_3774 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5332), .B(dp.rf._abc_6362_n5333), .Y(dp.rf._abc_6362_n4084) );
	NAND2X1 NAND2X1_3775 ( .gnd(gnd), .vdd(vdd), .A(dp.result_31_), .B(dp.rf._abc_6362_n5240), .Y(dp.rf._abc_6362_n5335) );
	NAND2X1 NAND2X1_3776 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_9_<31>), .B(dp.rf._abc_6362_n5242), .Y(dp.rf._abc_6362_n5336) );
	NAND2X1 NAND2X1_3777 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5335), .B(dp.rf._abc_6362_n5336), .Y(dp.rf._abc_6362_n4085) );
	INVX8 INVX8_37 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .Y(dp.rf._abc_6362_n5338) );
	NAND2X1 NAND2X1_3778 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<0>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5339) );
	INVX8 INVX8_38 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .Y(dp.rf._abc_6362_n5340) );
	INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<0>), .Y(dp.rf._abc_6362_n5341) );
	NOR2X1 NOR2X1_224 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5341), .Y(dp.rf._abc_6362_n5342) );
	NOR2X1 NOR2X1_225 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5342), .Y(dp.rf._abc_6362_n5343) );
	NAND2X1 NAND2X1_3779 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5339), .B(dp.rf._abc_6362_n5343), .Y(dp.rf._abc_6362_n5344) );
	NAND2X1 NAND2X1_3780 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<0>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5345) );
	INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<0>), .Y(dp.rf._abc_6362_n5346) );
	NOR2X1 NOR2X1_226 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5346), .Y(dp.rf._abc_6362_n5347) );
	NOR2X1 NOR2X1_227 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5347), .Y(dp.rf._abc_6362_n5348) );
	NAND2X1 NAND2X1_3781 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5345), .B(dp.rf._abc_6362_n5348), .Y(dp.rf._abc_6362_n5349) );
	NAND2X1 NAND2X1_3782 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5344), .B(dp.rf._abc_6362_n5349), .Y(dp.rf._abc_6362_n5350) );
	NAND2X1 NAND2X1_3783 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5350), .Y(dp.rf._abc_6362_n5351) );
	INVX8 INVX8_39 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .Y(dp.rf._abc_6362_n5352) );
	NAND2X1 NAND2X1_3784 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<0>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5353) );
	INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<0>), .Y(dp.rf._abc_6362_n5354) );
	NOR2X1 NOR2X1_228 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5354), .Y(dp.rf._abc_6362_n5355) );
	NOR2X1 NOR2X1_229 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5355), .Y(dp.rf._abc_6362_n5356) );
	NAND2X1 NAND2X1_3785 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5353), .B(dp.rf._abc_6362_n5356), .Y(dp.rf._abc_6362_n5357) );
	NAND2X1 NAND2X1_3786 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<0>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5358) );
	INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<0>), .Y(dp.rf._abc_6362_n5359) );
	NOR2X1 NOR2X1_230 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5359), .Y(dp.rf._abc_6362_n5360) );
	NOR2X1 NOR2X1_231 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5360), .Y(dp.rf._abc_6362_n5361) );
	NAND2X1 NAND2X1_3787 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5358), .B(dp.rf._abc_6362_n5361), .Y(dp.rf._abc_6362_n5362) );
	NAND2X1 NAND2X1_3788 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5357), .B(dp.rf._abc_6362_n5362), .Y(dp.rf._abc_6362_n5363) );
	NAND2X1 NAND2X1_3789 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5363), .Y(dp.rf._abc_6362_n5364) );
	NAND2X1 NAND2X1_3790 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5351), .B(dp.rf._abc_6362_n5364), .Y(dp.rf._abc_6362_n5365) );
	NOR2X1 NOR2X1_232 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5365), .Y(dp.rf._abc_6362_n5366) );
	INVX8 INVX8_40 ( .gnd(gnd), .vdd(vdd), .A(instr[25]), .Y(dp.rf._abc_6362_n5367) );
	NAND2X1 NAND2X1_3791 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<0>), .Y(dp.rf._abc_6362_n5368) );
	NAND2X1 NAND2X1_3792 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5368), .Y(dp.rf._abc_6362_n5369) );
	INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<0>), .Y(dp.rf._abc_6362_n5370) );
	NOR2X1 NOR2X1_233 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5370), .Y(dp.rf._abc_6362_n5371) );
	NOR2X1 NOR2X1_234 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5369), .B(dp.rf._abc_6362_n5371), .Y(dp.rf._abc_6362_n5372) );
	NAND2X1 NAND2X1_3793 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<0>), .Y(dp.rf._abc_6362_n5373) );
	NAND2X1 NAND2X1_3794 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5373), .Y(dp.rf._abc_6362_n5374) );
	INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<0>), .Y(dp.rf._abc_6362_n5375) );
	NOR2X1 NOR2X1_235 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5375), .Y(dp.rf._abc_6362_n5376) );
	NOR2X1 NOR2X1_236 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5374), .B(dp.rf._abc_6362_n5376), .Y(dp.rf._abc_6362_n5377) );
	OR2X2 OR2X2_30 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5372), .B(dp.rf._abc_6362_n5377), .Y(dp.rf._abc_6362_n5378) );
	NAND2X1 NAND2X1_3795 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5378), .Y(dp.rf._abc_6362_n5379) );
	NAND2X1 NAND2X1_3796 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<0>), .Y(dp.rf._abc_6362_n5380) );
	NAND2X1 NAND2X1_3797 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5380), .Y(dp.rf._abc_6362_n5381) );
	INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<0>), .Y(dp.rf._abc_6362_n5382) );
	NOR2X1 NOR2X1_237 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5382), .Y(dp.rf._abc_6362_n5383) );
	NOR2X1 NOR2X1_238 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5381), .B(dp.rf._abc_6362_n5383), .Y(dp.rf._abc_6362_n5384) );
	NAND2X1 NAND2X1_3798 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<0>), .Y(dp.rf._abc_6362_n5385) );
	NAND2X1 NAND2X1_3799 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5385), .Y(dp.rf._abc_6362_n5386) );
	INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<0>), .Y(dp.rf._abc_6362_n5387) );
	NOR2X1 NOR2X1_239 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5387), .Y(dp.rf._abc_6362_n5388) );
	NOR2X1 NOR2X1_240 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5386), .B(dp.rf._abc_6362_n5388), .Y(dp.rf._abc_6362_n5389) );
	OR2X2 OR2X2_31 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5384), .B(dp.rf._abc_6362_n5389), .Y(dp.rf._abc_6362_n5390) );
	NAND2X1 NAND2X1_3800 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5390), .Y(dp.rf._abc_6362_n5391) );
	AND2X2 AND2X2_76 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5391), .B(instr[24]), .Y(dp.rf._abc_6362_n5392) );
	NAND2X1 NAND2X1_3801 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5379), .B(dp.rf._abc_6362_n5392), .Y(dp.rf._abc_6362_n5393) );
	NAND2X1 NAND2X1_3802 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5393), .Y(dp.rf._abc_6362_n5394) );
	NOR2X1 NOR2X1_241 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5366), .B(dp.rf._abc_6362_n5394), .Y(dp.rf._abc_6362_n5395) );
	NOR2X1 NOR2X1_242 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(instr[22]), .Y(dp.rf._abc_6362_n5396) );
	INVX8 INVX8_41 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .Y(dp.rf._abc_6362_n5397) );
	NAND2X1 NAND2X1_3803 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n5398) );
	NOR2X1 NOR2X1_243 ( .gnd(gnd), .vdd(vdd), .A(instr[25]), .B(dp.rf._abc_6362_n5398), .Y(dp.rf._abc_6362_n5399) );
	NAND2X1 NAND2X1_3804 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5396), .B(dp.rf._abc_6362_n5399), .Y(dp.rf._abc_6362_n5400) );
	NAND2X1 NAND2X1_3805 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<0>), .Y(dp.rf._abc_6362_n5401) );
	NAND2X1 NAND2X1_3806 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5401), .Y(dp.rf._abc_6362_n5402) );
	INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<0>), .Y(dp.rf._abc_6362_n5403) );
	NOR2X1 NOR2X1_244 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5403), .Y(dp.rf._abc_6362_n5404) );
	NOR2X1 NOR2X1_245 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5402), .B(dp.rf._abc_6362_n5404), .Y(dp.rf._abc_6362_n5405) );
	NAND2X1 NAND2X1_3807 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<0>), .Y(dp.rf._abc_6362_n5406) );
	NAND2X1 NAND2X1_3808 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5406), .Y(dp.rf._abc_6362_n5407) );
	INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<0>), .Y(dp.rf._abc_6362_n5408) );
	NOR2X1 NOR2X1_246 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5408), .Y(dp.rf._abc_6362_n5409) );
	NOR2X1 NOR2X1_247 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5407), .B(dp.rf._abc_6362_n5409), .Y(dp.rf._abc_6362_n5410) );
	OR2X2 OR2X2_32 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5405), .B(dp.rf._abc_6362_n5410), .Y(dp.rf._abc_6362_n5411) );
	NAND2X1 NAND2X1_3809 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5411), .Y(dp.rf._abc_6362_n5412) );
	NAND2X1 NAND2X1_3810 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<0>), .Y(dp.rf._abc_6362_n5413) );
	NAND2X1 NAND2X1_3811 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5413), .Y(dp.rf._abc_6362_n5414) );
	INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<0>), .Y(dp.rf._abc_6362_n5415) );
	NOR2X1 NOR2X1_248 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5415), .Y(dp.rf._abc_6362_n5416) );
	NOR2X1 NOR2X1_249 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5414), .B(dp.rf._abc_6362_n5416), .Y(dp.rf._abc_6362_n5417) );
	NAND2X1 NAND2X1_3812 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<0>), .Y(dp.rf._abc_6362_n5418) );
	NAND2X1 NAND2X1_3813 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5418), .Y(dp.rf._abc_6362_n5419) );
	INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<0>), .Y(dp.rf._abc_6362_n5420) );
	NOR2X1 NOR2X1_250 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5420), .Y(dp.rf._abc_6362_n5421) );
	NOR2X1 NOR2X1_251 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5419), .B(dp.rf._abc_6362_n5421), .Y(dp.rf._abc_6362_n5422) );
	OR2X2 OR2X2_33 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5417), .B(dp.rf._abc_6362_n5422), .Y(dp.rf._abc_6362_n5423) );
	NAND2X1 NAND2X1_3814 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5423), .Y(dp.rf._abc_6362_n5424) );
	AND2X2 AND2X2_77 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5424), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n5425) );
	NAND2X1 NAND2X1_3815 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5412), .B(dp.rf._abc_6362_n5425), .Y(dp.rf._abc_6362_n5426) );
	NAND2X1 NAND2X1_3816 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<0>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5427) );
	NAND2X1 NAND2X1_3817 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<0>), .Y(dp.rf._abc_6362_n5428) );
	AND2X2 AND2X2_78 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5428), .B(instr[22]), .Y(dp.rf._abc_6362_n5429) );
	NAND2X1 NAND2X1_3818 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5427), .B(dp.rf._abc_6362_n5429), .Y(dp.rf._abc_6362_n5430) );
	NAND2X1 NAND2X1_3819 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<0>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5431) );
	NAND2X1 NAND2X1_3820 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<0>), .Y(dp.rf._abc_6362_n5432) );
	AND2X2 AND2X2_79 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5432), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5433) );
	NAND2X1 NAND2X1_3821 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5431), .B(dp.rf._abc_6362_n5433), .Y(dp.rf._abc_6362_n5434) );
	NAND2X1 NAND2X1_3822 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5430), .B(dp.rf._abc_6362_n5434), .Y(dp.rf._abc_6362_n5435) );
	AND2X2 AND2X2_80 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5435), .B(instr[23]), .Y(dp.rf._abc_6362_n5436) );
	NAND2X1 NAND2X1_3823 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<0>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5437) );
	NAND2X1 NAND2X1_3824 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<0>), .Y(dp.rf._abc_6362_n5438) );
	AND2X2 AND2X2_81 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5438), .B(instr[22]), .Y(dp.rf._abc_6362_n5439) );
	NAND2X1 NAND2X1_3825 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5437), .B(dp.rf._abc_6362_n5439), .Y(dp.rf._abc_6362_n5440) );
	NAND2X1 NAND2X1_3826 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<0>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5441) );
	NAND2X1 NAND2X1_3827 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<0>), .Y(dp.rf._abc_6362_n5442) );
	AND2X2 AND2X2_82 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5442), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5443) );
	NAND2X1 NAND2X1_3828 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5441), .B(dp.rf._abc_6362_n5443), .Y(dp.rf._abc_6362_n5444) );
	NAND2X1 NAND2X1_3829 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5440), .B(dp.rf._abc_6362_n5444), .Y(dp.rf._abc_6362_n5445) );
	NAND2X1 NAND2X1_3830 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5445), .Y(dp.rf._abc_6362_n5446) );
	NAND2X1 NAND2X1_3831 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5446), .Y(dp.rf._abc_6362_n5447) );
	NOR2X1 NOR2X1_252 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5436), .B(dp.rf._abc_6362_n5447), .Y(dp.rf._abc_6362_n5448) );
	NOR2X1 NOR2X1_253 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5448), .Y(dp.rf._abc_6362_n5449) );
	NAND2X1 NAND2X1_3832 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5426), .B(dp.rf._abc_6362_n5449), .Y(dp.rf._abc_6362_n5450) );
	NAND2X1 NAND2X1_3833 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n5450), .Y(dp.rf._abc_6362_n5451) );
	NOR2X1 NOR2X1_254 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5395), .B(dp.rf._abc_6362_n5451), .Y(dp.srca_0_) );
	NAND2X1 NAND2X1_3834 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<1>), .Y(dp.rf._abc_6362_n5453) );
	NAND2X1 NAND2X1_3835 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5453), .Y(dp.rf._abc_6362_n5454) );
	INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<1>), .Y(dp.rf._abc_6362_n5455) );
	NOR2X1 NOR2X1_255 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5455), .Y(dp.rf._abc_6362_n5456) );
	NOR2X1 NOR2X1_256 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5454), .B(dp.rf._abc_6362_n5456), .Y(dp.rf._abc_6362_n5457) );
	NAND2X1 NAND2X1_3836 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<1>), .Y(dp.rf._abc_6362_n5458) );
	NAND2X1 NAND2X1_3837 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5458), .Y(dp.rf._abc_6362_n5459) );
	INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<1>), .Y(dp.rf._abc_6362_n5460) );
	NOR2X1 NOR2X1_257 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5460), .Y(dp.rf._abc_6362_n5461) );
	NOR2X1 NOR2X1_258 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5459), .B(dp.rf._abc_6362_n5461), .Y(dp.rf._abc_6362_n5462) );
	NOR2X1 NOR2X1_259 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5457), .B(dp.rf._abc_6362_n5462), .Y(dp.rf._abc_6362_n5463) );
	NAND2X1 NAND2X1_3838 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5463), .Y(dp.rf._abc_6362_n5464) );
	NAND2X1 NAND2X1_3839 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<1>), .Y(dp.rf._abc_6362_n5465) );
	NAND2X1 NAND2X1_3840 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5465), .Y(dp.rf._abc_6362_n5466) );
	INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<1>), .Y(dp.rf._abc_6362_n5467) );
	NOR2X1 NOR2X1_260 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5467), .Y(dp.rf._abc_6362_n5468) );
	NOR2X1 NOR2X1_261 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5466), .B(dp.rf._abc_6362_n5468), .Y(dp.rf._abc_6362_n5469) );
	NAND2X1 NAND2X1_3841 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<1>), .Y(dp.rf._abc_6362_n5470) );
	NAND2X1 NAND2X1_3842 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5470), .Y(dp.rf._abc_6362_n5471) );
	INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<1>), .Y(dp.rf._abc_6362_n5472) );
	NOR2X1 NOR2X1_262 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5472), .Y(dp.rf._abc_6362_n5473) );
	NOR2X1 NOR2X1_263 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5471), .B(dp.rf._abc_6362_n5473), .Y(dp.rf._abc_6362_n5474) );
	NOR2X1 NOR2X1_264 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5469), .B(dp.rf._abc_6362_n5474), .Y(dp.rf._abc_6362_n5475) );
	NAND2X1 NAND2X1_3843 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5475), .Y(dp.rf._abc_6362_n5476) );
	NAND2X1 NAND2X1_3844 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5464), .B(dp.rf._abc_6362_n5476), .Y(dp.rf._abc_6362_n5477) );
	NAND2X1 NAND2X1_3845 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5477), .Y(dp.rf._abc_6362_n5478) );
	NAND2X1 NAND2X1_3846 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5478), .Y(dp.rf._abc_6362_n5479) );
	NAND2X1 NAND2X1_3847 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5480) );
	INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<1>), .Y(dp.rf._abc_6362_n5481) );
	NOR2X1 NOR2X1_265 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5481), .Y(dp.rf._abc_6362_n5482) );
	NOR2X1 NOR2X1_266 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5482), .Y(dp.rf._abc_6362_n5483) );
	NAND2X1 NAND2X1_3848 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5480), .B(dp.rf._abc_6362_n5483), .Y(dp.rf._abc_6362_n5484) );
	NAND2X1 NAND2X1_3849 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5485) );
	INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<1>), .Y(dp.rf._abc_6362_n5486) );
	NOR2X1 NOR2X1_267 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5486), .Y(dp.rf._abc_6362_n5487) );
	NOR2X1 NOR2X1_268 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5487), .Y(dp.rf._abc_6362_n5488) );
	NAND2X1 NAND2X1_3850 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5485), .B(dp.rf._abc_6362_n5488), .Y(dp.rf._abc_6362_n5489) );
	NAND2X1 NAND2X1_3851 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5484), .B(dp.rf._abc_6362_n5489), .Y(dp.rf._abc_6362_n5490) );
	NOR2X1 NOR2X1_269 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5490), .Y(dp.rf._abc_6362_n5491) );
	NAND2X1 NAND2X1_3852 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5492) );
	INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<1>), .Y(dp.rf._abc_6362_n5493) );
	NOR2X1 NOR2X1_270 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5493), .Y(dp.rf._abc_6362_n5494) );
	NOR2X1 NOR2X1_271 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5494), .Y(dp.rf._abc_6362_n5495) );
	NAND2X1 NAND2X1_3853 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5492), .B(dp.rf._abc_6362_n5495), .Y(dp.rf._abc_6362_n5496) );
	NAND2X1 NAND2X1_3854 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5497) );
	INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<1>), .Y(dp.rf._abc_6362_n5498) );
	NOR2X1 NOR2X1_272 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5498), .Y(dp.rf._abc_6362_n5499) );
	NOR2X1 NOR2X1_273 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5499), .Y(dp.rf._abc_6362_n5500) );
	NAND2X1 NAND2X1_3855 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5497), .B(dp.rf._abc_6362_n5500), .Y(dp.rf._abc_6362_n5501) );
	NAND2X1 NAND2X1_3856 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5496), .B(dp.rf._abc_6362_n5501), .Y(dp.rf._abc_6362_n5502) );
	NOR2X1 NOR2X1_274 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5502), .Y(dp.rf._abc_6362_n5503) );
	NOR2X1 NOR2X1_275 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5491), .B(dp.rf._abc_6362_n5503), .Y(dp.rf._abc_6362_n5504) );
	NOR2X1 NOR2X1_276 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5504), .Y(dp.rf._abc_6362_n5505) );
	NOR2X1 NOR2X1_277 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5479), .B(dp.rf._abc_6362_n5505), .Y(dp.rf._abc_6362_n5506) );
	NAND2X1 NAND2X1_3857 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<1>), .Y(dp.rf._abc_6362_n5507) );
	NAND2X1 NAND2X1_3858 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5508) );
	NAND2X1 NAND2X1_3859 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5507), .B(dp.rf._abc_6362_n5508), .Y(dp.rf._abc_6362_n5509) );
	NAND2X1 NAND2X1_3860 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5509), .Y(dp.rf._abc_6362_n5510) );
	NAND2X1 NAND2X1_3861 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<1>), .Y(dp.rf._abc_6362_n5511) );
	NAND2X1 NAND2X1_3862 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5512) );
	NAND2X1 NAND2X1_3863 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5511), .B(dp.rf._abc_6362_n5512), .Y(dp.rf._abc_6362_n5513) );
	NAND2X1 NAND2X1_3864 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5513), .Y(dp.rf._abc_6362_n5514) );
	AND2X2 AND2X2_83 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5510), .B(dp.rf._abc_6362_n5514), .Y(dp.rf._abc_6362_n5515) );
	NAND2X1 NAND2X1_3865 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5515), .Y(dp.rf._abc_6362_n5516) );
	NAND2X1 NAND2X1_3866 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<1>), .Y(dp.rf._abc_6362_n5517) );
	NAND2X1 NAND2X1_3867 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5518) );
	NAND2X1 NAND2X1_3868 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5517), .B(dp.rf._abc_6362_n5518), .Y(dp.rf._abc_6362_n5519) );
	NAND2X1 NAND2X1_3869 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5519), .Y(dp.rf._abc_6362_n5520) );
	NAND2X1 NAND2X1_3870 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<1>), .Y(dp.rf._abc_6362_n5521) );
	NAND2X1 NAND2X1_3871 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5522) );
	NAND2X1 NAND2X1_3872 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5521), .B(dp.rf._abc_6362_n5522), .Y(dp.rf._abc_6362_n5523) );
	NAND2X1 NAND2X1_3873 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5523), .Y(dp.rf._abc_6362_n5524) );
	AND2X2 AND2X2_84 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5520), .B(dp.rf._abc_6362_n5524), .Y(dp.rf._abc_6362_n5525) );
	NAND2X1 NAND2X1_3874 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5525), .Y(dp.rf._abc_6362_n5526) );
	AND2X2 AND2X2_85 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5526), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n5527) );
	NAND2X1 NAND2X1_3875 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5516), .B(dp.rf._abc_6362_n5527), .Y(dp.rf._abc_6362_n5528) );
	NAND2X1 NAND2X1_3876 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5529) );
	NAND2X1 NAND2X1_3877 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<1>), .Y(dp.rf._abc_6362_n5530) );
	AND2X2 AND2X2_86 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5530), .B(instr[22]), .Y(dp.rf._abc_6362_n5531) );
	NAND2X1 NAND2X1_3878 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5529), .B(dp.rf._abc_6362_n5531), .Y(dp.rf._abc_6362_n5532) );
	NAND2X1 NAND2X1_3879 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5533) );
	NAND2X1 NAND2X1_3880 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<1>), .Y(dp.rf._abc_6362_n5534) );
	AND2X2 AND2X2_87 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5534), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5535) );
	NAND2X1 NAND2X1_3881 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5533), .B(dp.rf._abc_6362_n5535), .Y(dp.rf._abc_6362_n5536) );
	NAND2X1 NAND2X1_3882 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5532), .B(dp.rf._abc_6362_n5536), .Y(dp.rf._abc_6362_n5537) );
	AND2X2 AND2X2_88 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5537), .B(instr[23]), .Y(dp.rf._abc_6362_n5538) );
	NAND2X1 NAND2X1_3883 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5539) );
	NAND2X1 NAND2X1_3884 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<1>), .Y(dp.rf._abc_6362_n5540) );
	AND2X2 AND2X2_89 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5540), .B(instr[22]), .Y(dp.rf._abc_6362_n5541) );
	NAND2X1 NAND2X1_3885 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5539), .B(dp.rf._abc_6362_n5541), .Y(dp.rf._abc_6362_n5542) );
	NAND2X1 NAND2X1_3886 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<1>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5543) );
	NAND2X1 NAND2X1_3887 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<1>), .Y(dp.rf._abc_6362_n5544) );
	AND2X2 AND2X2_90 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5544), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5545) );
	NAND2X1 NAND2X1_3888 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5543), .B(dp.rf._abc_6362_n5545), .Y(dp.rf._abc_6362_n5546) );
	NAND2X1 NAND2X1_3889 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5542), .B(dp.rf._abc_6362_n5546), .Y(dp.rf._abc_6362_n5547) );
	NAND2X1 NAND2X1_3890 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5547), .Y(dp.rf._abc_6362_n5548) );
	NAND2X1 NAND2X1_3891 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5548), .Y(dp.rf._abc_6362_n5549) );
	NOR2X1 NOR2X1_278 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5538), .B(dp.rf._abc_6362_n5549), .Y(dp.rf._abc_6362_n5550) );
	NOR2X1 NOR2X1_279 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5550), .Y(dp.rf._abc_6362_n5551) );
	NAND2X1 NAND2X1_3892 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5528), .B(dp.rf._abc_6362_n5551), .Y(dp.rf._abc_6362_n5552) );
	NAND2X1 NAND2X1_3893 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n5552), .Y(dp.rf._abc_6362_n5553) );
	NOR2X1 NOR2X1_280 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5506), .B(dp.rf._abc_6362_n5553), .Y(dp.srca_1_) );
	NAND2X1 NAND2X1_3894 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<2>), .Y(dp.rf._abc_6362_n5555) );
	NAND2X1 NAND2X1_3895 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5555), .Y(dp.rf._abc_6362_n5556) );
	INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<2>), .Y(dp.rf._abc_6362_n5557) );
	NOR2X1 NOR2X1_281 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5557), .Y(dp.rf._abc_6362_n5558) );
	NOR2X1 NOR2X1_282 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5556), .B(dp.rf._abc_6362_n5558), .Y(dp.rf._abc_6362_n5559) );
	NAND2X1 NAND2X1_3896 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<2>), .Y(dp.rf._abc_6362_n5560) );
	NAND2X1 NAND2X1_3897 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5560), .Y(dp.rf._abc_6362_n5561) );
	INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<2>), .Y(dp.rf._abc_6362_n5562) );
	NOR2X1 NOR2X1_283 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5562), .Y(dp.rf._abc_6362_n5563) );
	NOR2X1 NOR2X1_284 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5561), .B(dp.rf._abc_6362_n5563), .Y(dp.rf._abc_6362_n5564) );
	NOR2X1 NOR2X1_285 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5559), .B(dp.rf._abc_6362_n5564), .Y(dp.rf._abc_6362_n5565) );
	NAND2X1 NAND2X1_3898 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5565), .Y(dp.rf._abc_6362_n5566) );
	NAND2X1 NAND2X1_3899 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<2>), .Y(dp.rf._abc_6362_n5567) );
	NAND2X1 NAND2X1_3900 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5567), .Y(dp.rf._abc_6362_n5568) );
	INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<2>), .Y(dp.rf._abc_6362_n5569) );
	NOR2X1 NOR2X1_286 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5569), .Y(dp.rf._abc_6362_n5570) );
	NOR2X1 NOR2X1_287 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5568), .B(dp.rf._abc_6362_n5570), .Y(dp.rf._abc_6362_n5571) );
	NAND2X1 NAND2X1_3901 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<2>), .Y(dp.rf._abc_6362_n5572) );
	NAND2X1 NAND2X1_3902 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5572), .Y(dp.rf._abc_6362_n5573) );
	INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<2>), .Y(dp.rf._abc_6362_n5574) );
	NOR2X1 NOR2X1_288 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5574), .Y(dp.rf._abc_6362_n5575) );
	NOR2X1 NOR2X1_289 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5573), .B(dp.rf._abc_6362_n5575), .Y(dp.rf._abc_6362_n5576) );
	NOR2X1 NOR2X1_290 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5571), .B(dp.rf._abc_6362_n5576), .Y(dp.rf._abc_6362_n5577) );
	NAND2X1 NAND2X1_3903 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5577), .Y(dp.rf._abc_6362_n5578) );
	NAND2X1 NAND2X1_3904 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5566), .B(dp.rf._abc_6362_n5578), .Y(dp.rf._abc_6362_n5579) );
	NAND2X1 NAND2X1_3905 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5579), .Y(dp.rf._abc_6362_n5580) );
	NAND2X1 NAND2X1_3906 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5580), .Y(dp.rf._abc_6362_n5581) );
	NAND2X1 NAND2X1_3907 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5582) );
	INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<2>), .Y(dp.rf._abc_6362_n5583) );
	NOR2X1 NOR2X1_291 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5583), .Y(dp.rf._abc_6362_n5584) );
	NOR2X1 NOR2X1_292 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5584), .Y(dp.rf._abc_6362_n5585) );
	NAND2X1 NAND2X1_3908 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5582), .B(dp.rf._abc_6362_n5585), .Y(dp.rf._abc_6362_n5586) );
	NAND2X1 NAND2X1_3909 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5587) );
	INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<2>), .Y(dp.rf._abc_6362_n5588) );
	NOR2X1 NOR2X1_293 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5588), .Y(dp.rf._abc_6362_n5589) );
	NOR2X1 NOR2X1_294 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5589), .Y(dp.rf._abc_6362_n5590) );
	NAND2X1 NAND2X1_3910 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5587), .B(dp.rf._abc_6362_n5590), .Y(dp.rf._abc_6362_n5591) );
	NAND2X1 NAND2X1_3911 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5586), .B(dp.rf._abc_6362_n5591), .Y(dp.rf._abc_6362_n5592) );
	NOR2X1 NOR2X1_295 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5592), .Y(dp.rf._abc_6362_n5593) );
	NAND2X1 NAND2X1_3912 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5594) );
	INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<2>), .Y(dp.rf._abc_6362_n5595) );
	NOR2X1 NOR2X1_296 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5595), .Y(dp.rf._abc_6362_n5596) );
	NOR2X1 NOR2X1_297 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5596), .Y(dp.rf._abc_6362_n5597) );
	NAND2X1 NAND2X1_3913 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5594), .B(dp.rf._abc_6362_n5597), .Y(dp.rf._abc_6362_n5598) );
	NAND2X1 NAND2X1_3914 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5599) );
	INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<2>), .Y(dp.rf._abc_6362_n5600) );
	NOR2X1 NOR2X1_298 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5600), .Y(dp.rf._abc_6362_n5601) );
	NOR2X1 NOR2X1_299 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5601), .Y(dp.rf._abc_6362_n5602) );
	NAND2X1 NAND2X1_3915 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5599), .B(dp.rf._abc_6362_n5602), .Y(dp.rf._abc_6362_n5603) );
	NAND2X1 NAND2X1_3916 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5598), .B(dp.rf._abc_6362_n5603), .Y(dp.rf._abc_6362_n5604) );
	NOR2X1 NOR2X1_300 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5604), .Y(dp.rf._abc_6362_n5605) );
	NOR2X1 NOR2X1_301 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5593), .B(dp.rf._abc_6362_n5605), .Y(dp.rf._abc_6362_n5606) );
	NOR2X1 NOR2X1_302 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5606), .Y(dp.rf._abc_6362_n5607) );
	NOR2X1 NOR2X1_303 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5581), .B(dp.rf._abc_6362_n5607), .Y(dp.rf._abc_6362_n5608) );
	NAND2X1 NAND2X1_3917 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<2>), .Y(dp.rf._abc_6362_n5609) );
	NAND2X1 NAND2X1_3918 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5610) );
	NAND2X1 NAND2X1_3919 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5609), .B(dp.rf._abc_6362_n5610), .Y(dp.rf._abc_6362_n5611) );
	NAND2X1 NAND2X1_3920 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5611), .Y(dp.rf._abc_6362_n5612) );
	NAND2X1 NAND2X1_3921 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<2>), .Y(dp.rf._abc_6362_n5613) );
	NAND2X1 NAND2X1_3922 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5614) );
	NAND2X1 NAND2X1_3923 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5613), .B(dp.rf._abc_6362_n5614), .Y(dp.rf._abc_6362_n5615) );
	NAND2X1 NAND2X1_3924 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5615), .Y(dp.rf._abc_6362_n5616) );
	AND2X2 AND2X2_91 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5612), .B(dp.rf._abc_6362_n5616), .Y(dp.rf._abc_6362_n5617) );
	NAND2X1 NAND2X1_3925 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5617), .Y(dp.rf._abc_6362_n5618) );
	NAND2X1 NAND2X1_3926 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<2>), .Y(dp.rf._abc_6362_n5619) );
	NAND2X1 NAND2X1_3927 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5620) );
	NAND2X1 NAND2X1_3928 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5619), .B(dp.rf._abc_6362_n5620), .Y(dp.rf._abc_6362_n5621) );
	NAND2X1 NAND2X1_3929 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5621), .Y(dp.rf._abc_6362_n5622) );
	NAND2X1 NAND2X1_3930 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<2>), .Y(dp.rf._abc_6362_n5623) );
	NAND2X1 NAND2X1_3931 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5624) );
	NAND2X1 NAND2X1_3932 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5623), .B(dp.rf._abc_6362_n5624), .Y(dp.rf._abc_6362_n5625) );
	NAND2X1 NAND2X1_3933 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5625), .Y(dp.rf._abc_6362_n5626) );
	AND2X2 AND2X2_92 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5622), .B(dp.rf._abc_6362_n5626), .Y(dp.rf._abc_6362_n5627) );
	NAND2X1 NAND2X1_3934 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5627), .Y(dp.rf._abc_6362_n5628) );
	AND2X2 AND2X2_93 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5628), .B(instr[24]), .Y(dp.rf._abc_6362_n5629) );
	NAND2X1 NAND2X1_3935 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5618), .B(dp.rf._abc_6362_n5629), .Y(dp.rf._abc_6362_n5630) );
	NAND2X1 NAND2X1_3936 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5631) );
	NAND2X1 NAND2X1_3937 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<2>), .Y(dp.rf._abc_6362_n5632) );
	AND2X2 AND2X2_94 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5632), .B(instr[22]), .Y(dp.rf._abc_6362_n5633) );
	NAND2X1 NAND2X1_3938 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5631), .B(dp.rf._abc_6362_n5633), .Y(dp.rf._abc_6362_n5634) );
	NAND2X1 NAND2X1_3939 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5635) );
	NAND2X1 NAND2X1_3940 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<2>), .Y(dp.rf._abc_6362_n5636) );
	AND2X2 AND2X2_95 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5636), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5637) );
	NAND2X1 NAND2X1_3941 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5635), .B(dp.rf._abc_6362_n5637), .Y(dp.rf._abc_6362_n5638) );
	NAND2X1 NAND2X1_3942 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5634), .B(dp.rf._abc_6362_n5638), .Y(dp.rf._abc_6362_n5639) );
	AND2X2 AND2X2_96 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5639), .B(instr[23]), .Y(dp.rf._abc_6362_n5640) );
	NAND2X1 NAND2X1_3943 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5641) );
	NAND2X1 NAND2X1_3944 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<2>), .Y(dp.rf._abc_6362_n5642) );
	AND2X2 AND2X2_97 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5642), .B(instr[22]), .Y(dp.rf._abc_6362_n5643) );
	NAND2X1 NAND2X1_3945 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5641), .B(dp.rf._abc_6362_n5643), .Y(dp.rf._abc_6362_n5644) );
	NAND2X1 NAND2X1_3946 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<2>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5645) );
	NAND2X1 NAND2X1_3947 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<2>), .Y(dp.rf._abc_6362_n5646) );
	AND2X2 AND2X2_98 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5646), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5647) );
	NAND2X1 NAND2X1_3948 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5645), .B(dp.rf._abc_6362_n5647), .Y(dp.rf._abc_6362_n5648) );
	NAND2X1 NAND2X1_3949 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5644), .B(dp.rf._abc_6362_n5648), .Y(dp.rf._abc_6362_n5649) );
	NAND2X1 NAND2X1_3950 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5649), .Y(dp.rf._abc_6362_n5650) );
	NAND2X1 NAND2X1_3951 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n5650), .Y(dp.rf._abc_6362_n5651) );
	NOR2X1 NOR2X1_304 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5640), .B(dp.rf._abc_6362_n5651), .Y(dp.rf._abc_6362_n5652) );
	NOR2X1 NOR2X1_305 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5652), .Y(dp.rf._abc_6362_n5653) );
	NAND2X1 NAND2X1_3952 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5630), .B(dp.rf._abc_6362_n5653), .Y(dp.rf._abc_6362_n5654) );
	NAND2X1 NAND2X1_3953 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n5654), .Y(dp.rf._abc_6362_n5655) );
	NOR2X1 NOR2X1_306 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5608), .B(dp.rf._abc_6362_n5655), .Y(dp.srca_2_) );
	NAND2X1 NAND2X1_3954 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<3>), .Y(dp.rf._abc_6362_n5657) );
	NAND2X1 NAND2X1_3955 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5657), .Y(dp.rf._abc_6362_n5658) );
	INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<3>), .Y(dp.rf._abc_6362_n5659) );
	NOR2X1 NOR2X1_307 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5659), .Y(dp.rf._abc_6362_n5660) );
	NOR2X1 NOR2X1_308 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5658), .B(dp.rf._abc_6362_n5660), .Y(dp.rf._abc_6362_n5661) );
	NAND2X1 NAND2X1_3956 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<3>), .Y(dp.rf._abc_6362_n5662) );
	NAND2X1 NAND2X1_3957 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5662), .Y(dp.rf._abc_6362_n5663) );
	INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<3>), .Y(dp.rf._abc_6362_n5664) );
	NOR2X1 NOR2X1_309 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5664), .Y(dp.rf._abc_6362_n5665) );
	NOR2X1 NOR2X1_310 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5663), .B(dp.rf._abc_6362_n5665), .Y(dp.rf._abc_6362_n5666) );
	NOR2X1 NOR2X1_311 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5661), .B(dp.rf._abc_6362_n5666), .Y(dp.rf._abc_6362_n5667) );
	NAND2X1 NAND2X1_3958 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5667), .Y(dp.rf._abc_6362_n5668) );
	NAND2X1 NAND2X1_3959 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<3>), .Y(dp.rf._abc_6362_n5669) );
	NAND2X1 NAND2X1_3960 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5669), .Y(dp.rf._abc_6362_n5670) );
	INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<3>), .Y(dp.rf._abc_6362_n5671) );
	NOR2X1 NOR2X1_312 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5671), .Y(dp.rf._abc_6362_n5672) );
	NOR2X1 NOR2X1_313 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5670), .B(dp.rf._abc_6362_n5672), .Y(dp.rf._abc_6362_n5673) );
	NAND2X1 NAND2X1_3961 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<3>), .Y(dp.rf._abc_6362_n5674) );
	NAND2X1 NAND2X1_3962 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5674), .Y(dp.rf._abc_6362_n5675) );
	INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<3>), .Y(dp.rf._abc_6362_n5676) );
	NOR2X1 NOR2X1_314 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5676), .Y(dp.rf._abc_6362_n5677) );
	NOR2X1 NOR2X1_315 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5675), .B(dp.rf._abc_6362_n5677), .Y(dp.rf._abc_6362_n5678) );
	NOR2X1 NOR2X1_316 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5673), .B(dp.rf._abc_6362_n5678), .Y(dp.rf._abc_6362_n5679) );
	NAND2X1 NAND2X1_3963 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5679), .Y(dp.rf._abc_6362_n5680) );
	NAND2X1 NAND2X1_3964 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5668), .B(dp.rf._abc_6362_n5680), .Y(dp.rf._abc_6362_n5681) );
	NAND2X1 NAND2X1_3965 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5681), .Y(dp.rf._abc_6362_n5682) );
	NAND2X1 NAND2X1_3966 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5682), .Y(dp.rf._abc_6362_n5683) );
	NAND2X1 NAND2X1_3967 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5684) );
	INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<3>), .Y(dp.rf._abc_6362_n5685) );
	NOR2X1 NOR2X1_317 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5685), .Y(dp.rf._abc_6362_n5686) );
	NOR2X1 NOR2X1_318 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5686), .Y(dp.rf._abc_6362_n5687) );
	NAND2X1 NAND2X1_3968 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5684), .B(dp.rf._abc_6362_n5687), .Y(dp.rf._abc_6362_n5688) );
	NAND2X1 NAND2X1_3969 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5689) );
	INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<3>), .Y(dp.rf._abc_6362_n5690) );
	NOR2X1 NOR2X1_319 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5690), .Y(dp.rf._abc_6362_n5691) );
	NOR2X1 NOR2X1_320 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5691), .Y(dp.rf._abc_6362_n5692) );
	NAND2X1 NAND2X1_3970 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5689), .B(dp.rf._abc_6362_n5692), .Y(dp.rf._abc_6362_n5693) );
	NAND2X1 NAND2X1_3971 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5688), .B(dp.rf._abc_6362_n5693), .Y(dp.rf._abc_6362_n5694) );
	NOR2X1 NOR2X1_321 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5694), .Y(dp.rf._abc_6362_n5695) );
	NAND2X1 NAND2X1_3972 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5696) );
	INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<3>), .Y(dp.rf._abc_6362_n5697) );
	NOR2X1 NOR2X1_322 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5697), .Y(dp.rf._abc_6362_n5698) );
	NOR2X1 NOR2X1_323 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5698), .Y(dp.rf._abc_6362_n5699) );
	NAND2X1 NAND2X1_3973 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5696), .B(dp.rf._abc_6362_n5699), .Y(dp.rf._abc_6362_n5700) );
	NAND2X1 NAND2X1_3974 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5701) );
	INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<3>), .Y(dp.rf._abc_6362_n5702) );
	NOR2X1 NOR2X1_324 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n5702), .Y(dp.rf._abc_6362_n5703) );
	NOR2X1 NOR2X1_325 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5703), .Y(dp.rf._abc_6362_n5704) );
	NAND2X1 NAND2X1_3975 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5701), .B(dp.rf._abc_6362_n5704), .Y(dp.rf._abc_6362_n5705) );
	NAND2X1 NAND2X1_3976 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5700), .B(dp.rf._abc_6362_n5705), .Y(dp.rf._abc_6362_n5706) );
	NOR2X1 NOR2X1_326 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5706), .Y(dp.rf._abc_6362_n5707) );
	NOR2X1 NOR2X1_327 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5695), .B(dp.rf._abc_6362_n5707), .Y(dp.rf._abc_6362_n5708) );
	NOR2X1 NOR2X1_328 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5708), .Y(dp.rf._abc_6362_n5709) );
	NOR2X1 NOR2X1_329 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5683), .B(dp.rf._abc_6362_n5709), .Y(dp.rf._abc_6362_n5710) );
	NAND2X1 NAND2X1_3977 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<3>), .Y(dp.rf._abc_6362_n5711) );
	NAND2X1 NAND2X1_3978 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5712) );
	NAND2X1 NAND2X1_3979 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5711), .B(dp.rf._abc_6362_n5712), .Y(dp.rf._abc_6362_n5713) );
	NAND2X1 NAND2X1_3980 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5713), .Y(dp.rf._abc_6362_n5714) );
	NAND2X1 NAND2X1_3981 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<3>), .Y(dp.rf._abc_6362_n5715) );
	NAND2X1 NAND2X1_3982 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5716) );
	NAND2X1 NAND2X1_3983 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5715), .B(dp.rf._abc_6362_n5716), .Y(dp.rf._abc_6362_n5717) );
	NAND2X1 NAND2X1_3984 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5717), .Y(dp.rf._abc_6362_n5718) );
	AND2X2 AND2X2_99 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5714), .B(dp.rf._abc_6362_n5718), .Y(dp.rf._abc_6362_n5719) );
	NAND2X1 NAND2X1_3985 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5719), .Y(dp.rf._abc_6362_n5720) );
	NAND2X1 NAND2X1_3986 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<3>), .Y(dp.rf._abc_6362_n5721) );
	NAND2X1 NAND2X1_3987 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5722) );
	NAND2X1 NAND2X1_3988 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5721), .B(dp.rf._abc_6362_n5722), .Y(dp.rf._abc_6362_n5723) );
	NAND2X1 NAND2X1_3989 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5723), .Y(dp.rf._abc_6362_n5724) );
	NAND2X1 NAND2X1_3990 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<3>), .Y(dp.rf._abc_6362_n5725) );
	NAND2X1 NAND2X1_3991 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5726) );
	NAND2X1 NAND2X1_3992 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5725), .B(dp.rf._abc_6362_n5726), .Y(dp.rf._abc_6362_n5727) );
	NAND2X1 NAND2X1_3993 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5727), .Y(dp.rf._abc_6362_n5728) );
	AND2X2 AND2X2_100 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5724), .B(dp.rf._abc_6362_n5728), .Y(dp.rf._abc_6362_n5729) );
	NAND2X1 NAND2X1_3994 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5729), .Y(dp.rf._abc_6362_n5730) );
	AND2X2 AND2X2_101 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5730), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n5731) );
	NAND2X1 NAND2X1_3995 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5720), .B(dp.rf._abc_6362_n5731), .Y(dp.rf._abc_6362_n5732) );
	NAND2X1 NAND2X1_3996 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5733) );
	NAND2X1 NAND2X1_3997 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<3>), .Y(dp.rf._abc_6362_n5734) );
	AND2X2 AND2X2_102 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5734), .B(instr[22]), .Y(dp.rf._abc_6362_n5735) );
	NAND2X1 NAND2X1_3998 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5733), .B(dp.rf._abc_6362_n5735), .Y(dp.rf._abc_6362_n5736) );
	NAND2X1 NAND2X1_3999 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5737) );
	NAND2X1 NAND2X1_4000 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<3>), .Y(dp.rf._abc_6362_n5738) );
	AND2X2 AND2X2_103 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5738), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5739) );
	NAND2X1 NAND2X1_4001 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5737), .B(dp.rf._abc_6362_n5739), .Y(dp.rf._abc_6362_n5740) );
	NAND2X1 NAND2X1_4002 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5736), .B(dp.rf._abc_6362_n5740), .Y(dp.rf._abc_6362_n5741) );
	AND2X2 AND2X2_104 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5741), .B(instr[23]), .Y(dp.rf._abc_6362_n5742) );
	NAND2X1 NAND2X1_4003 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5743) );
	NAND2X1 NAND2X1_4004 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<3>), .Y(dp.rf._abc_6362_n5744) );
	AND2X2 AND2X2_105 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5744), .B(instr[22]), .Y(dp.rf._abc_6362_n5745) );
	NAND2X1 NAND2X1_4005 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5743), .B(dp.rf._abc_6362_n5745), .Y(dp.rf._abc_6362_n5746) );
	NAND2X1 NAND2X1_4006 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<3>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5747) );
	NAND2X1 NAND2X1_4007 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<3>), .Y(dp.rf._abc_6362_n5748) );
	AND2X2 AND2X2_106 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5748), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5749) );
	NAND2X1 NAND2X1_4008 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5747), .B(dp.rf._abc_6362_n5749), .Y(dp.rf._abc_6362_n5750) );
	NAND2X1 NAND2X1_4009 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5746), .B(dp.rf._abc_6362_n5750), .Y(dp.rf._abc_6362_n5751) );
	NAND2X1 NAND2X1_4010 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5751), .Y(dp.rf._abc_6362_n5752) );
	NAND2X1 NAND2X1_4011 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5752), .Y(dp.rf._abc_6362_n5753) );
	NOR2X1 NOR2X1_330 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5742), .B(dp.rf._abc_6362_n5753), .Y(dp.rf._abc_6362_n5754) );
	NOR2X1 NOR2X1_331 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5754), .Y(dp.rf._abc_6362_n5755) );
	NAND2X1 NAND2X1_4012 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5732), .B(dp.rf._abc_6362_n5755), .Y(dp.rf._abc_6362_n5756) );
	NAND2X1 NAND2X1_4013 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n5756), .Y(dp.rf._abc_6362_n5757) );
	NOR2X1 NOR2X1_332 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5710), .B(dp.rf._abc_6362_n5757), .Y(dp.srca_3_) );
	NAND2X1 NAND2X1_4014 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<4>), .Y(dp.rf._abc_6362_n5759) );
	NAND2X1 NAND2X1_4015 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5760) );
	NAND2X1 NAND2X1_4016 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5759), .B(dp.rf._abc_6362_n5760), .Y(dp.rf._abc_6362_n5761) );
	NAND2X1 NAND2X1_4017 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5761), .Y(dp.rf._abc_6362_n5762) );
	NAND2X1 NAND2X1_4018 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<4>), .Y(dp.rf._abc_6362_n5763) );
	NAND2X1 NAND2X1_4019 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5764) );
	NAND2X1 NAND2X1_4020 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5763), .B(dp.rf._abc_6362_n5764), .Y(dp.rf._abc_6362_n5765) );
	NAND2X1 NAND2X1_4021 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5765), .Y(dp.rf._abc_6362_n5766) );
	NAND2X1 NAND2X1_4022 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5762), .B(dp.rf._abc_6362_n5766), .Y(dp.rf._abc_6362_n5767) );
	NOR2X1 NOR2X1_333 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5767), .Y(dp.rf._abc_6362_n5768) );
	NAND2X1 NAND2X1_4023 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<4>), .Y(dp.rf._abc_6362_n5769) );
	NAND2X1 NAND2X1_4024 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5770) );
	NAND2X1 NAND2X1_4025 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5769), .B(dp.rf._abc_6362_n5770), .Y(dp.rf._abc_6362_n5771) );
	NAND2X1 NAND2X1_4026 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5771), .Y(dp.rf._abc_6362_n5772) );
	NAND2X1 NAND2X1_4027 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<4>), .Y(dp.rf._abc_6362_n5773) );
	NAND2X1 NAND2X1_4028 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5774) );
	NAND2X1 NAND2X1_4029 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5773), .B(dp.rf._abc_6362_n5774), .Y(dp.rf._abc_6362_n5775) );
	NAND2X1 NAND2X1_4030 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5775), .Y(dp.rf._abc_6362_n5776) );
	AND2X2 AND2X2_107 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5772), .B(dp.rf._abc_6362_n5776), .Y(dp.rf._abc_6362_n5777) );
	NAND2X1 NAND2X1_4031 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5777), .Y(dp.rf._abc_6362_n5778) );
	NAND2X1 NAND2X1_4032 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n5778), .Y(dp.rf._abc_6362_n5779) );
	NOR2X1 NOR2X1_334 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5768), .B(dp.rf._abc_6362_n5779), .Y(dp.rf._abc_6362_n5780) );
	NAND2X1 NAND2X1_4033 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<4>), .Y(dp.rf._abc_6362_n5781) );
	NAND2X1 NAND2X1_4034 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5781), .Y(dp.rf._abc_6362_n5782) );
	INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<4>), .Y(dp.rf._abc_6362_n5783) );
	NOR2X1 NOR2X1_335 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5783), .Y(dp.rf._abc_6362_n5784) );
	NOR2X1 NOR2X1_336 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5782), .B(dp.rf._abc_6362_n5784), .Y(dp.rf._abc_6362_n5785) );
	NAND2X1 NAND2X1_4035 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<4>), .Y(dp.rf._abc_6362_n5786) );
	NAND2X1 NAND2X1_4036 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5786), .Y(dp.rf._abc_6362_n5787) );
	INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<4>), .Y(dp.rf._abc_6362_n5788) );
	NOR2X1 NOR2X1_337 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5788), .Y(dp.rf._abc_6362_n5789) );
	NOR2X1 NOR2X1_338 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5787), .B(dp.rf._abc_6362_n5789), .Y(dp.rf._abc_6362_n5790) );
	NOR2X1 NOR2X1_339 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5785), .B(dp.rf._abc_6362_n5790), .Y(dp.rf._abc_6362_n5791) );
	NAND2X1 NAND2X1_4037 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5791), .Y(dp.rf._abc_6362_n5792) );
	NAND2X1 NAND2X1_4038 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<4>), .Y(dp.rf._abc_6362_n5793) );
	NAND2X1 NAND2X1_4039 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5793), .Y(dp.rf._abc_6362_n5794) );
	INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<4>), .Y(dp.rf._abc_6362_n5795) );
	NOR2X1 NOR2X1_340 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5795), .Y(dp.rf._abc_6362_n5796) );
	NOR2X1 NOR2X1_341 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5794), .B(dp.rf._abc_6362_n5796), .Y(dp.rf._abc_6362_n5797) );
	NAND2X1 NAND2X1_4040 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<4>), .Y(dp.rf._abc_6362_n5798) );
	NAND2X1 NAND2X1_4041 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5798), .Y(dp.rf._abc_6362_n5799) );
	INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<4>), .Y(dp.rf._abc_6362_n5800) );
	NOR2X1 NOR2X1_342 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5800), .Y(dp.rf._abc_6362_n5801) );
	NOR2X1 NOR2X1_343 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5799), .B(dp.rf._abc_6362_n5801), .Y(dp.rf._abc_6362_n5802) );
	NOR2X1 NOR2X1_344 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5797), .B(dp.rf._abc_6362_n5802), .Y(dp.rf._abc_6362_n5803) );
	NAND2X1 NAND2X1_4042 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5803), .Y(dp.rf._abc_6362_n5804) );
	NAND2X1 NAND2X1_4043 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5792), .B(dp.rf._abc_6362_n5804), .Y(dp.rf._abc_6362_n5805) );
	NAND2X1 NAND2X1_4044 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5805), .Y(dp.rf._abc_6362_n5806) );
	NAND2X1 NAND2X1_4045 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5806), .Y(dp.rf._abc_6362_n5807) );
	NOR2X1 NOR2X1_345 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5780), .B(dp.rf._abc_6362_n5807), .Y(dp.rf._abc_6362_n5808) );
	NAND2X1 NAND2X1_4046 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<4>), .Y(dp.rf._abc_6362_n5809) );
	NAND2X1 NAND2X1_4047 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5810) );
	NAND2X1 NAND2X1_4048 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5809), .B(dp.rf._abc_6362_n5810), .Y(dp.rf._abc_6362_n5811) );
	NAND2X1 NAND2X1_4049 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5811), .Y(dp.rf._abc_6362_n5812) );
	NAND2X1 NAND2X1_4050 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<4>), .Y(dp.rf._abc_6362_n5813) );
	NAND2X1 NAND2X1_4051 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5814) );
	NAND2X1 NAND2X1_4052 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5813), .B(dp.rf._abc_6362_n5814), .Y(dp.rf._abc_6362_n5815) );
	NAND2X1 NAND2X1_4053 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5815), .Y(dp.rf._abc_6362_n5816) );
	AND2X2 AND2X2_108 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5812), .B(dp.rf._abc_6362_n5816), .Y(dp.rf._abc_6362_n5817) );
	NAND2X1 NAND2X1_4054 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5817), .Y(dp.rf._abc_6362_n5818) );
	NAND2X1 NAND2X1_4055 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<4>), .Y(dp.rf._abc_6362_n5819) );
	NAND2X1 NAND2X1_4056 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5820) );
	NAND2X1 NAND2X1_4057 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5819), .B(dp.rf._abc_6362_n5820), .Y(dp.rf._abc_6362_n5821) );
	NAND2X1 NAND2X1_4058 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5821), .Y(dp.rf._abc_6362_n5822) );
	NAND2X1 NAND2X1_4059 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<4>), .Y(dp.rf._abc_6362_n5823) );
	NAND2X1 NAND2X1_4060 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5824) );
	NAND2X1 NAND2X1_4061 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5823), .B(dp.rf._abc_6362_n5824), .Y(dp.rf._abc_6362_n5825) );
	NAND2X1 NAND2X1_4062 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5825), .Y(dp.rf._abc_6362_n5826) );
	AND2X2 AND2X2_109 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5822), .B(dp.rf._abc_6362_n5826), .Y(dp.rf._abc_6362_n5827) );
	NAND2X1 NAND2X1_4063 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5827), .Y(dp.rf._abc_6362_n5828) );
	AND2X2 AND2X2_110 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5828), .B(instr[24]), .Y(dp.rf._abc_6362_n5829) );
	NAND2X1 NAND2X1_4064 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5818), .B(dp.rf._abc_6362_n5829), .Y(dp.rf._abc_6362_n5830) );
	NAND2X1 NAND2X1_4065 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5831) );
	NAND2X1 NAND2X1_4066 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<4>), .Y(dp.rf._abc_6362_n5832) );
	AND2X2 AND2X2_111 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5832), .B(instr[22]), .Y(dp.rf._abc_6362_n5833) );
	NAND2X1 NAND2X1_4067 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5831), .B(dp.rf._abc_6362_n5833), .Y(dp.rf._abc_6362_n5834) );
	NAND2X1 NAND2X1_4068 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5835) );
	NAND2X1 NAND2X1_4069 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<4>), .Y(dp.rf._abc_6362_n5836) );
	AND2X2 AND2X2_112 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5836), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5837) );
	NAND2X1 NAND2X1_4070 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5835), .B(dp.rf._abc_6362_n5837), .Y(dp.rf._abc_6362_n5838) );
	NAND2X1 NAND2X1_4071 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5834), .B(dp.rf._abc_6362_n5838), .Y(dp.rf._abc_6362_n5839) );
	AND2X2 AND2X2_113 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5839), .B(instr[23]), .Y(dp.rf._abc_6362_n5840) );
	NAND2X1 NAND2X1_4072 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5841) );
	NAND2X1 NAND2X1_4073 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<4>), .Y(dp.rf._abc_6362_n5842) );
	AND2X2 AND2X2_114 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5842), .B(instr[22]), .Y(dp.rf._abc_6362_n5843) );
	NAND2X1 NAND2X1_4074 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5841), .B(dp.rf._abc_6362_n5843), .Y(dp.rf._abc_6362_n5844) );
	NAND2X1 NAND2X1_4075 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<4>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5845) );
	NAND2X1 NAND2X1_4076 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<4>), .Y(dp.rf._abc_6362_n5846) );
	AND2X2 AND2X2_115 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5846), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5847) );
	NAND2X1 NAND2X1_4077 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5845), .B(dp.rf._abc_6362_n5847), .Y(dp.rf._abc_6362_n5848) );
	NAND2X1 NAND2X1_4078 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5844), .B(dp.rf._abc_6362_n5848), .Y(dp.rf._abc_6362_n5849) );
	NAND2X1 NAND2X1_4079 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5849), .Y(dp.rf._abc_6362_n5850) );
	NAND2X1 NAND2X1_4080 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n5850), .Y(dp.rf._abc_6362_n5851) );
	NOR2X1 NOR2X1_346 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5840), .B(dp.rf._abc_6362_n5851), .Y(dp.rf._abc_6362_n5852) );
	NOR2X1 NOR2X1_347 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5852), .Y(dp.rf._abc_6362_n5853) );
	NAND2X1 NAND2X1_4081 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5830), .B(dp.rf._abc_6362_n5853), .Y(dp.rf._abc_6362_n5854) );
	NAND2X1 NAND2X1_4082 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n5854), .Y(dp.rf._abc_6362_n5855) );
	NOR2X1 NOR2X1_348 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5808), .B(dp.rf._abc_6362_n5855), .Y(dp.srca_4_) );
	NAND2X1 NAND2X1_4083 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<5>), .Y(dp.rf._abc_6362_n5857) );
	NAND2X1 NAND2X1_4084 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<5>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5858) );
	NAND2X1 NAND2X1_4085 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5857), .B(dp.rf._abc_6362_n5858), .Y(dp.rf._abc_6362_n5859) );
	NAND2X1 NAND2X1_4086 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5859), .Y(dp.rf._abc_6362_n5860) );
	NAND2X1 NAND2X1_4087 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<5>), .Y(dp.rf._abc_6362_n5861) );
	NAND2X1 NAND2X1_4088 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<5>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5862) );
	NAND2X1 NAND2X1_4089 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5861), .B(dp.rf._abc_6362_n5862), .Y(dp.rf._abc_6362_n5863) );
	NAND2X1 NAND2X1_4090 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5863), .Y(dp.rf._abc_6362_n5864) );
	NAND2X1 NAND2X1_4091 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5860), .B(dp.rf._abc_6362_n5864), .Y(dp.rf._abc_6362_n5865) );
	NOR2X1 NOR2X1_349 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5865), .Y(dp.rf._abc_6362_n5866) );
	NAND2X1 NAND2X1_4092 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<5>), .Y(dp.rf._abc_6362_n5867) );
	NAND2X1 NAND2X1_4093 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<5>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5868) );
	NAND2X1 NAND2X1_4094 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5867), .B(dp.rf._abc_6362_n5868), .Y(dp.rf._abc_6362_n5869) );
	NAND2X1 NAND2X1_4095 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5869), .Y(dp.rf._abc_6362_n5870) );
	NAND2X1 NAND2X1_4096 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<5>), .Y(dp.rf._abc_6362_n5871) );
	NAND2X1 NAND2X1_4097 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<5>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5872) );
	NAND2X1 NAND2X1_4098 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5871), .B(dp.rf._abc_6362_n5872), .Y(dp.rf._abc_6362_n5873) );
	NAND2X1 NAND2X1_4099 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5873), .Y(dp.rf._abc_6362_n5874) );
	AND2X2 AND2X2_116 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5870), .B(dp.rf._abc_6362_n5874), .Y(dp.rf._abc_6362_n5875) );
	NAND2X1 NAND2X1_4100 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5875), .Y(dp.rf._abc_6362_n5876) );
	NAND2X1 NAND2X1_4101 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5876), .Y(dp.rf._abc_6362_n5877) );
	NOR2X1 NOR2X1_350 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5866), .B(dp.rf._abc_6362_n5877), .Y(dp.rf._abc_6362_n5878) );
	NAND2X1 NAND2X1_4102 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<5>), .Y(dp.rf._abc_6362_n5879) );
	NAND2X1 NAND2X1_4103 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<5>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5880) );
	NAND2X1 NAND2X1_4104 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5879), .B(dp.rf._abc_6362_n5880), .Y(dp.rf._abc_6362_n5881) );
	NAND2X1 NAND2X1_4105 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5881), .Y(dp.rf._abc_6362_n5882) );
	NAND2X1 NAND2X1_4106 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<5>), .Y(dp.rf._abc_6362_n5883) );
	NAND2X1 NAND2X1_4107 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<5>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5884) );
	NAND2X1 NAND2X1_4108 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5883), .B(dp.rf._abc_6362_n5884), .Y(dp.rf._abc_6362_n5885) );
	NAND2X1 NAND2X1_4109 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5885), .Y(dp.rf._abc_6362_n5886) );
	AND2X2 AND2X2_117 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5882), .B(dp.rf._abc_6362_n5886), .Y(dp.rf._abc_6362_n5887) );
	NAND2X1 NAND2X1_4110 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5887), .Y(dp.rf._abc_6362_n5888) );
	NAND2X1 NAND2X1_4111 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<5>), .Y(dp.rf._abc_6362_n5889) );
	NAND2X1 NAND2X1_4112 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5889), .Y(dp.rf._abc_6362_n5890) );
	AND2X2 AND2X2_118 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf.rf_2_<5>), .Y(dp.rf._abc_6362_n5891) );
	NOR2X1 NOR2X1_351 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5890), .B(dp.rf._abc_6362_n5891), .Y(dp.rf._abc_6362_n5892) );
	NAND2X1 NAND2X1_4113 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<5>), .Y(dp.rf._abc_6362_n5893) );
	NAND2X1 NAND2X1_4114 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5893), .Y(dp.rf._abc_6362_n5894) );
	INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<5>), .Y(dp.rf._abc_6362_n5895) );
	NOR2X1 NOR2X1_352 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5895), .Y(dp.rf._abc_6362_n5896) );
	NOR2X1 NOR2X1_353 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5894), .B(dp.rf._abc_6362_n5896), .Y(dp.rf._abc_6362_n5897) );
	OR2X2 OR2X2_34 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5892), .B(dp.rf._abc_6362_n5897), .Y(dp.rf._abc_6362_n5898) );
	NAND2X1 NAND2X1_4115 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5898), .Y(dp.rf._abc_6362_n5899) );
	AND2X2 AND2X2_119 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5899), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n5900) );
	NAND2X1 NAND2X1_4116 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5888), .B(dp.rf._abc_6362_n5900), .Y(dp.rf._abc_6362_n5901) );
	NAND2X1 NAND2X1_4117 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5901), .Y(dp.rf._abc_6362_n5902) );
	NOR2X1 NOR2X1_354 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5878), .B(dp.rf._abc_6362_n5902), .Y(dp.rf._abc_6362_n5903) );
	NAND2X1 NAND2X1_4118 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<5>), .Y(dp.rf._abc_6362_n5904) );
	NAND2X1 NAND2X1_4119 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5904), .Y(dp.rf._abc_6362_n5905) );
	INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<5>), .Y(dp.rf._abc_6362_n5906) );
	NOR2X1 NOR2X1_355 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5906), .Y(dp.rf._abc_6362_n5907) );
	NOR2X1 NOR2X1_356 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5905), .B(dp.rf._abc_6362_n5907), .Y(dp.rf._abc_6362_n5908) );
	NAND2X1 NAND2X1_4120 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<5>), .Y(dp.rf._abc_6362_n5909) );
	NAND2X1 NAND2X1_4121 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5909), .Y(dp.rf._abc_6362_n5910) );
	INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<5>), .Y(dp.rf._abc_6362_n5911) );
	NOR2X1 NOR2X1_357 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5911), .Y(dp.rf._abc_6362_n5912) );
	NOR2X1 NOR2X1_358 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5910), .B(dp.rf._abc_6362_n5912), .Y(dp.rf._abc_6362_n5913) );
	OR2X2 OR2X2_35 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5908), .B(dp.rf._abc_6362_n5913), .Y(dp.rf._abc_6362_n5914) );
	NAND2X1 NAND2X1_4122 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5914), .Y(dp.rf._abc_6362_n5915) );
	NAND2X1 NAND2X1_4123 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<5>), .Y(dp.rf._abc_6362_n5916) );
	NAND2X1 NAND2X1_4124 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5916), .Y(dp.rf._abc_6362_n5917) );
	INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<5>), .Y(dp.rf._abc_6362_n5918) );
	NOR2X1 NOR2X1_359 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5918), .Y(dp.rf._abc_6362_n5919) );
	NOR2X1 NOR2X1_360 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5917), .B(dp.rf._abc_6362_n5919), .Y(dp.rf._abc_6362_n5920) );
	NAND2X1 NAND2X1_4125 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<5>), .Y(dp.rf._abc_6362_n5921) );
	NAND2X1 NAND2X1_4126 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5921), .Y(dp.rf._abc_6362_n5922) );
	INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<5>), .Y(dp.rf._abc_6362_n5923) );
	NOR2X1 NOR2X1_361 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n5923), .Y(dp.rf._abc_6362_n5924) );
	NOR2X1 NOR2X1_362 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5922), .B(dp.rf._abc_6362_n5924), .Y(dp.rf._abc_6362_n5925) );
	OR2X2 OR2X2_36 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5920), .B(dp.rf._abc_6362_n5925), .Y(dp.rf._abc_6362_n5926) );
	NAND2X1 NAND2X1_4127 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5926), .Y(dp.rf._abc_6362_n5927) );
	AND2X2 AND2X2_120 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5927), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n5928) );
	NAND2X1 NAND2X1_4128 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5915), .B(dp.rf._abc_6362_n5928), .Y(dp.rf._abc_6362_n5929) );
	NAND2X1 NAND2X1_4129 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<5>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5930) );
	NAND2X1 NAND2X1_4130 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<5>), .Y(dp.rf._abc_6362_n5931) );
	AND2X2 AND2X2_121 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5931), .B(instr[22]), .Y(dp.rf._abc_6362_n5932) );
	NAND2X1 NAND2X1_4131 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5930), .B(dp.rf._abc_6362_n5932), .Y(dp.rf._abc_6362_n5933) );
	NAND2X1 NAND2X1_4132 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<5>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5934) );
	NAND2X1 NAND2X1_4133 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<5>), .Y(dp.rf._abc_6362_n5935) );
	AND2X2 AND2X2_122 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5935), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5936) );
	NAND2X1 NAND2X1_4134 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5934), .B(dp.rf._abc_6362_n5936), .Y(dp.rf._abc_6362_n5937) );
	NAND2X1 NAND2X1_4135 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5933), .B(dp.rf._abc_6362_n5937), .Y(dp.rf._abc_6362_n5938) );
	AND2X2 AND2X2_123 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5938), .B(instr[23]), .Y(dp.rf._abc_6362_n5939) );
	NAND2X1 NAND2X1_4136 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<5>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5940) );
	NAND2X1 NAND2X1_4137 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<5>), .Y(dp.rf._abc_6362_n5941) );
	AND2X2 AND2X2_124 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5941), .B(instr[22]), .Y(dp.rf._abc_6362_n5942) );
	NAND2X1 NAND2X1_4138 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5940), .B(dp.rf._abc_6362_n5942), .Y(dp.rf._abc_6362_n5943) );
	NAND2X1 NAND2X1_4139 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<5>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5944) );
	NAND2X1 NAND2X1_4140 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<5>), .Y(dp.rf._abc_6362_n5945) );
	AND2X2 AND2X2_125 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5945), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n5946) );
	NAND2X1 NAND2X1_4141 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5944), .B(dp.rf._abc_6362_n5946), .Y(dp.rf._abc_6362_n5947) );
	NAND2X1 NAND2X1_4142 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5943), .B(dp.rf._abc_6362_n5947), .Y(dp.rf._abc_6362_n5948) );
	NAND2X1 NAND2X1_4143 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5948), .Y(dp.rf._abc_6362_n5949) );
	NAND2X1 NAND2X1_4144 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5949), .Y(dp.rf._abc_6362_n5950) );
	NOR2X1 NOR2X1_363 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5939), .B(dp.rf._abc_6362_n5950), .Y(dp.rf._abc_6362_n5951) );
	NOR2X1 NOR2X1_364 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5951), .Y(dp.rf._abc_6362_n5952) );
	NAND2X1 NAND2X1_4145 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5929), .B(dp.rf._abc_6362_n5952), .Y(dp.rf._abc_6362_n5953) );
	NAND2X1 NAND2X1_4146 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n5953), .Y(dp.rf._abc_6362_n5954) );
	NOR2X1 NOR2X1_365 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5903), .B(dp.rf._abc_6362_n5954), .Y(dp.srca_5_) );
	NAND2X1 NAND2X1_4147 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<6>), .Y(dp.rf._abc_6362_n5956) );
	NAND2X1 NAND2X1_4148 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5957) );
	NAND2X1 NAND2X1_4149 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5956), .B(dp.rf._abc_6362_n5957), .Y(dp.rf._abc_6362_n5958) );
	NAND2X1 NAND2X1_4150 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5958), .Y(dp.rf._abc_6362_n5959) );
	NAND2X1 NAND2X1_4151 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<6>), .Y(dp.rf._abc_6362_n5960) );
	NAND2X1 NAND2X1_4152 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5961) );
	NAND2X1 NAND2X1_4153 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5960), .B(dp.rf._abc_6362_n5961), .Y(dp.rf._abc_6362_n5962) );
	NAND2X1 NAND2X1_4154 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5962), .Y(dp.rf._abc_6362_n5963) );
	NAND2X1 NAND2X1_4155 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5959), .B(dp.rf._abc_6362_n5963), .Y(dp.rf._abc_6362_n5964) );
	NOR2X1 NOR2X1_366 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5964), .Y(dp.rf._abc_6362_n5965) );
	NAND2X1 NAND2X1_4156 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<6>), .Y(dp.rf._abc_6362_n5966) );
	NAND2X1 NAND2X1_4157 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5967) );
	NAND2X1 NAND2X1_4158 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5966), .B(dp.rf._abc_6362_n5967), .Y(dp.rf._abc_6362_n5968) );
	NAND2X1 NAND2X1_4159 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5968), .Y(dp.rf._abc_6362_n5969) );
	NAND2X1 NAND2X1_4160 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<6>), .Y(dp.rf._abc_6362_n5970) );
	NAND2X1 NAND2X1_4161 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5971) );
	NAND2X1 NAND2X1_4162 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5970), .B(dp.rf._abc_6362_n5971), .Y(dp.rf._abc_6362_n5972) );
	NAND2X1 NAND2X1_4163 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5972), .Y(dp.rf._abc_6362_n5973) );
	AND2X2 AND2X2_126 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5969), .B(dp.rf._abc_6362_n5973), .Y(dp.rf._abc_6362_n5974) );
	NAND2X1 NAND2X1_4164 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5974), .Y(dp.rf._abc_6362_n5975) );
	NAND2X1 NAND2X1_4165 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n5975), .Y(dp.rf._abc_6362_n5976) );
	NOR2X1 NOR2X1_367 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5965), .B(dp.rf._abc_6362_n5976), .Y(dp.rf._abc_6362_n5977) );
	NAND2X1 NAND2X1_4166 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<6>), .Y(dp.rf._abc_6362_n5978) );
	NAND2X1 NAND2X1_4167 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5979) );
	NAND2X1 NAND2X1_4168 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5978), .B(dp.rf._abc_6362_n5979), .Y(dp.rf._abc_6362_n5980) );
	NAND2X1 NAND2X1_4169 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5980), .Y(dp.rf._abc_6362_n5981) );
	NAND2X1 NAND2X1_4170 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<6>), .Y(dp.rf._abc_6362_n5982) );
	NAND2X1 NAND2X1_4171 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5983) );
	NAND2X1 NAND2X1_4172 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5982), .B(dp.rf._abc_6362_n5983), .Y(dp.rf._abc_6362_n5984) );
	NAND2X1 NAND2X1_4173 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5984), .Y(dp.rf._abc_6362_n5985) );
	NAND2X1 NAND2X1_4174 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5981), .B(dp.rf._abc_6362_n5985), .Y(dp.rf._abc_6362_n5986) );
	NAND2X1 NAND2X1_4175 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n5986), .Y(dp.rf._abc_6362_n5987) );
	NAND2X1 NAND2X1_4176 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<6>), .Y(dp.rf._abc_6362_n5988) );
	NAND2X1 NAND2X1_4177 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5989) );
	NAND2X1 NAND2X1_4178 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5988), .B(dp.rf._abc_6362_n5989), .Y(dp.rf._abc_6362_n5990) );
	NAND2X1 NAND2X1_4179 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n5990), .Y(dp.rf._abc_6362_n5991) );
	NAND2X1 NAND2X1_4180 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<6>), .Y(dp.rf._abc_6362_n5992) );
	NAND2X1 NAND2X1_4181 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n5993) );
	NAND2X1 NAND2X1_4182 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5992), .B(dp.rf._abc_6362_n5993), .Y(dp.rf._abc_6362_n5994) );
	NAND2X1 NAND2X1_4183 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n5994), .Y(dp.rf._abc_6362_n5995) );
	NAND2X1 NAND2X1_4184 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5991), .B(dp.rf._abc_6362_n5995), .Y(dp.rf._abc_6362_n5996) );
	NAND2X1 NAND2X1_4185 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n5996), .Y(dp.rf._abc_6362_n5997) );
	NAND2X1 NAND2X1_4186 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5987), .B(dp.rf._abc_6362_n5997), .Y(dp.rf._abc_6362_n5998) );
	NAND2X1 NAND2X1_4187 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n5998), .Y(dp.rf._abc_6362_n5999) );
	NAND2X1 NAND2X1_4188 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n5999), .Y(dp.rf._abc_6362_n6000) );
	NOR2X1 NOR2X1_368 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5977), .B(dp.rf._abc_6362_n6000), .Y(dp.rf._abc_6362_n6001) );
	NAND2X1 NAND2X1_4189 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<6>), .Y(dp.rf._abc_6362_n6002) );
	NAND2X1 NAND2X1_4190 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6002), .Y(dp.rf._abc_6362_n6003) );
	INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<6>), .Y(dp.rf._abc_6362_n6004) );
	NOR2X1 NOR2X1_369 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6004), .Y(dp.rf._abc_6362_n6005) );
	NOR2X1 NOR2X1_370 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6003), .B(dp.rf._abc_6362_n6005), .Y(dp.rf._abc_6362_n6006) );
	NAND2X1 NAND2X1_4191 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<6>), .Y(dp.rf._abc_6362_n6007) );
	NAND2X1 NAND2X1_4192 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6007), .Y(dp.rf._abc_6362_n6008) );
	INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<6>), .Y(dp.rf._abc_6362_n6009) );
	NOR2X1 NOR2X1_371 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6009), .Y(dp.rf._abc_6362_n6010) );
	NOR2X1 NOR2X1_372 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6008), .B(dp.rf._abc_6362_n6010), .Y(dp.rf._abc_6362_n6011) );
	OR2X2 OR2X2_37 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6006), .B(dp.rf._abc_6362_n6011), .Y(dp.rf._abc_6362_n6012) );
	NAND2X1 NAND2X1_4193 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6012), .Y(dp.rf._abc_6362_n6013) );
	NAND2X1 NAND2X1_4194 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<6>), .Y(dp.rf._abc_6362_n6014) );
	NAND2X1 NAND2X1_4195 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6014), .Y(dp.rf._abc_6362_n6015) );
	INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<6>), .Y(dp.rf._abc_6362_n6016) );
	NOR2X1 NOR2X1_373 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6016), .Y(dp.rf._abc_6362_n6017) );
	NOR2X1 NOR2X1_374 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6015), .B(dp.rf._abc_6362_n6017), .Y(dp.rf._abc_6362_n6018) );
	NAND2X1 NAND2X1_4196 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<6>), .Y(dp.rf._abc_6362_n6019) );
	NAND2X1 NAND2X1_4197 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6019), .Y(dp.rf._abc_6362_n6020) );
	INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<6>), .Y(dp.rf._abc_6362_n6021) );
	NOR2X1 NOR2X1_375 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6021), .Y(dp.rf._abc_6362_n6022) );
	NOR2X1 NOR2X1_376 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6020), .B(dp.rf._abc_6362_n6022), .Y(dp.rf._abc_6362_n6023) );
	OR2X2 OR2X2_38 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6018), .B(dp.rf._abc_6362_n6023), .Y(dp.rf._abc_6362_n6024) );
	NAND2X1 NAND2X1_4198 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6024), .Y(dp.rf._abc_6362_n6025) );
	AND2X2 AND2X2_127 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6025), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n6026) );
	NAND2X1 NAND2X1_4199 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6013), .B(dp.rf._abc_6362_n6026), .Y(dp.rf._abc_6362_n6027) );
	NAND2X1 NAND2X1_4200 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6028) );
	NAND2X1 NAND2X1_4201 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<6>), .Y(dp.rf._abc_6362_n6029) );
	AND2X2 AND2X2_128 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6029), .B(instr[22]), .Y(dp.rf._abc_6362_n6030) );
	NAND2X1 NAND2X1_4202 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6028), .B(dp.rf._abc_6362_n6030), .Y(dp.rf._abc_6362_n6031) );
	NAND2X1 NAND2X1_4203 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6032) );
	NAND2X1 NAND2X1_4204 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<6>), .Y(dp.rf._abc_6362_n6033) );
	AND2X2 AND2X2_129 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6033), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6034) );
	NAND2X1 NAND2X1_4205 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6032), .B(dp.rf._abc_6362_n6034), .Y(dp.rf._abc_6362_n6035) );
	NAND2X1 NAND2X1_4206 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6031), .B(dp.rf._abc_6362_n6035), .Y(dp.rf._abc_6362_n6036) );
	AND2X2 AND2X2_130 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6036), .B(instr[23]), .Y(dp.rf._abc_6362_n6037) );
	NAND2X1 NAND2X1_4207 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6038) );
	NAND2X1 NAND2X1_4208 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<6>), .Y(dp.rf._abc_6362_n6039) );
	AND2X2 AND2X2_131 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6039), .B(instr[22]), .Y(dp.rf._abc_6362_n6040) );
	NAND2X1 NAND2X1_4209 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6038), .B(dp.rf._abc_6362_n6040), .Y(dp.rf._abc_6362_n6041) );
	NAND2X1 NAND2X1_4210 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<6>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6042) );
	NAND2X1 NAND2X1_4211 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<6>), .Y(dp.rf._abc_6362_n6043) );
	AND2X2 AND2X2_132 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6043), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6044) );
	NAND2X1 NAND2X1_4212 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6042), .B(dp.rf._abc_6362_n6044), .Y(dp.rf._abc_6362_n6045) );
	NAND2X1 NAND2X1_4213 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6041), .B(dp.rf._abc_6362_n6045), .Y(dp.rf._abc_6362_n6046) );
	NAND2X1 NAND2X1_4214 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6046), .Y(dp.rf._abc_6362_n6047) );
	NAND2X1 NAND2X1_4215 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6047), .Y(dp.rf._abc_6362_n6048) );
	NOR2X1 NOR2X1_377 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6037), .B(dp.rf._abc_6362_n6048), .Y(dp.rf._abc_6362_n6049) );
	NOR2X1 NOR2X1_378 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6049), .Y(dp.rf._abc_6362_n6050) );
	NAND2X1 NAND2X1_4216 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6027), .B(dp.rf._abc_6362_n6050), .Y(dp.rf._abc_6362_n6051) );
	NAND2X1 NAND2X1_4217 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n6051), .Y(dp.rf._abc_6362_n6052) );
	NOR2X1 NOR2X1_379 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6001), .B(dp.rf._abc_6362_n6052), .Y(dp.srca_6_) );
	NAND2X1 NAND2X1_4218 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<7>), .Y(dp.rf._abc_6362_n6054) );
	NAND2X1 NAND2X1_4219 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6054), .Y(dp.rf._abc_6362_n6055) );
	INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<7>), .Y(dp.rf._abc_6362_n6056) );
	NOR2X1 NOR2X1_380 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6056), .Y(dp.rf._abc_6362_n6057) );
	NOR2X1 NOR2X1_381 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6055), .B(dp.rf._abc_6362_n6057), .Y(dp.rf._abc_6362_n6058) );
	NAND2X1 NAND2X1_4220 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<7>), .Y(dp.rf._abc_6362_n6059) );
	NAND2X1 NAND2X1_4221 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6059), .Y(dp.rf._abc_6362_n6060) );
	INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<7>), .Y(dp.rf._abc_6362_n6061) );
	NOR2X1 NOR2X1_382 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6061), .Y(dp.rf._abc_6362_n6062) );
	NOR2X1 NOR2X1_383 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6060), .B(dp.rf._abc_6362_n6062), .Y(dp.rf._abc_6362_n6063) );
	NOR2X1 NOR2X1_384 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6058), .B(dp.rf._abc_6362_n6063), .Y(dp.rf._abc_6362_n6064) );
	NAND2X1 NAND2X1_4222 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6064), .Y(dp.rf._abc_6362_n6065) );
	NAND2X1 NAND2X1_4223 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<7>), .Y(dp.rf._abc_6362_n6066) );
	NAND2X1 NAND2X1_4224 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6066), .Y(dp.rf._abc_6362_n6067) );
	INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<7>), .Y(dp.rf._abc_6362_n6068) );
	NOR2X1 NOR2X1_385 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6068), .Y(dp.rf._abc_6362_n6069) );
	NOR2X1 NOR2X1_386 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6067), .B(dp.rf._abc_6362_n6069), .Y(dp.rf._abc_6362_n6070) );
	NAND2X1 NAND2X1_4225 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<7>), .Y(dp.rf._abc_6362_n6071) );
	NAND2X1 NAND2X1_4226 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6071), .Y(dp.rf._abc_6362_n6072) );
	INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<7>), .Y(dp.rf._abc_6362_n6073) );
	NOR2X1 NOR2X1_387 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6073), .Y(dp.rf._abc_6362_n6074) );
	NOR2X1 NOR2X1_388 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6072), .B(dp.rf._abc_6362_n6074), .Y(dp.rf._abc_6362_n6075) );
	NOR2X1 NOR2X1_389 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6070), .B(dp.rf._abc_6362_n6075), .Y(dp.rf._abc_6362_n6076) );
	NAND2X1 NAND2X1_4227 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6076), .Y(dp.rf._abc_6362_n6077) );
	NAND2X1 NAND2X1_4228 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6065), .B(dp.rf._abc_6362_n6077), .Y(dp.rf._abc_6362_n6078) );
	NAND2X1 NAND2X1_4229 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6078), .Y(dp.rf._abc_6362_n6079) );
	NAND2X1 NAND2X1_4230 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<7>), .Y(dp.rf._abc_6362_n6080) );
	NAND2X1 NAND2X1_4231 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<7>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6081) );
	NAND2X1 NAND2X1_4232 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6080), .B(dp.rf._abc_6362_n6081), .Y(dp.rf._abc_6362_n6082) );
	NAND2X1 NAND2X1_4233 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6082), .Y(dp.rf._abc_6362_n6083) );
	NAND2X1 NAND2X1_4234 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<7>), .Y(dp.rf._abc_6362_n6084) );
	NAND2X1 NAND2X1_4235 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<7>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6085) );
	NAND2X1 NAND2X1_4236 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6084), .B(dp.rf._abc_6362_n6085), .Y(dp.rf._abc_6362_n6086) );
	NAND2X1 NAND2X1_4237 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6086), .Y(dp.rf._abc_6362_n6087) );
	AND2X2 AND2X2_133 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6083), .B(dp.rf._abc_6362_n6087), .Y(dp.rf._abc_6362_n6088) );
	NAND2X1 NAND2X1_4238 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6088), .Y(dp.rf._abc_6362_n6089) );
	NAND2X1 NAND2X1_4239 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<7>), .Y(dp.rf._abc_6362_n6090) );
	NAND2X1 NAND2X1_4240 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6090), .Y(dp.rf._abc_6362_n6091) );
	AND2X2 AND2X2_134 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf.rf_2_<7>), .Y(dp.rf._abc_6362_n6092) );
	NOR2X1 NOR2X1_390 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6091), .B(dp.rf._abc_6362_n6092), .Y(dp.rf._abc_6362_n6093) );
	NAND2X1 NAND2X1_4241 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<7>), .Y(dp.rf._abc_6362_n6094) );
	NAND2X1 NAND2X1_4242 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6094), .Y(dp.rf._abc_6362_n6095) );
	INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<7>), .Y(dp.rf._abc_6362_n6096) );
	NOR2X1 NOR2X1_391 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6096), .Y(dp.rf._abc_6362_n6097) );
	NOR2X1 NOR2X1_392 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6095), .B(dp.rf._abc_6362_n6097), .Y(dp.rf._abc_6362_n6098) );
	OR2X2 OR2X2_39 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6093), .B(dp.rf._abc_6362_n6098), .Y(dp.rf._abc_6362_n6099) );
	NAND2X1 NAND2X1_4243 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6099), .Y(dp.rf._abc_6362_n6100) );
	AND2X2 AND2X2_135 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6100), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n6101) );
	NAND2X1 NAND2X1_4244 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6089), .B(dp.rf._abc_6362_n6101), .Y(dp.rf._abc_6362_n6102) );
	NAND2X1 NAND2X1_4245 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6079), .B(dp.rf._abc_6362_n6102), .Y(dp.rf._abc_6362_n6103) );
	NOR2X1 NOR2X1_393 ( .gnd(gnd), .vdd(vdd), .A(instr[25]), .B(dp.rf._abc_6362_n6103), .Y(dp.rf._abc_6362_n6104) );
	NAND2X1 NAND2X1_4246 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<7>), .Y(dp.rf._abc_6362_n6105) );
	NAND2X1 NAND2X1_4247 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6105), .Y(dp.rf._abc_6362_n6106) );
	INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<7>), .Y(dp.rf._abc_6362_n6107) );
	NOR2X1 NOR2X1_394 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6107), .Y(dp.rf._abc_6362_n6108) );
	NOR2X1 NOR2X1_395 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6106), .B(dp.rf._abc_6362_n6108), .Y(dp.rf._abc_6362_n6109) );
	NAND2X1 NAND2X1_4248 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<7>), .Y(dp.rf._abc_6362_n6110) );
	NAND2X1 NAND2X1_4249 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6110), .Y(dp.rf._abc_6362_n6111) );
	INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<7>), .Y(dp.rf._abc_6362_n6112) );
	NOR2X1 NOR2X1_396 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6112), .Y(dp.rf._abc_6362_n6113) );
	NOR2X1 NOR2X1_397 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6111), .B(dp.rf._abc_6362_n6113), .Y(dp.rf._abc_6362_n6114) );
	OR2X2 OR2X2_40 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6109), .B(dp.rf._abc_6362_n6114), .Y(dp.rf._abc_6362_n6115) );
	NAND2X1 NAND2X1_4250 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6115), .Y(dp.rf._abc_6362_n6116) );
	NAND2X1 NAND2X1_4251 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<7>), .Y(dp.rf._abc_6362_n6117) );
	NAND2X1 NAND2X1_4252 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6117), .Y(dp.rf._abc_6362_n6118) );
	INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<7>), .Y(dp.rf._abc_6362_n6119) );
	NOR2X1 NOR2X1_398 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6119), .Y(dp.rf._abc_6362_n6120) );
	NOR2X1 NOR2X1_399 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6118), .B(dp.rf._abc_6362_n6120), .Y(dp.rf._abc_6362_n6121) );
	NAND2X1 NAND2X1_4253 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<7>), .Y(dp.rf._abc_6362_n6122) );
	NAND2X1 NAND2X1_4254 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6122), .Y(dp.rf._abc_6362_n6123) );
	INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<7>), .Y(dp.rf._abc_6362_n6124) );
	NOR2X1 NOR2X1_400 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6124), .Y(dp.rf._abc_6362_n6125) );
	NOR2X1 NOR2X1_401 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6123), .B(dp.rf._abc_6362_n6125), .Y(dp.rf._abc_6362_n6126) );
	OR2X2 OR2X2_41 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6121), .B(dp.rf._abc_6362_n6126), .Y(dp.rf._abc_6362_n6127) );
	NAND2X1 NAND2X1_4255 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6127), .Y(dp.rf._abc_6362_n6128) );
	AND2X2 AND2X2_136 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6128), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n6129) );
	NAND2X1 NAND2X1_4256 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6116), .B(dp.rf._abc_6362_n6129), .Y(dp.rf._abc_6362_n6130) );
	NAND2X1 NAND2X1_4257 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<7>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6131) );
	NAND2X1 NAND2X1_4258 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<7>), .Y(dp.rf._abc_6362_n6132) );
	AND2X2 AND2X2_137 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6132), .B(instr[22]), .Y(dp.rf._abc_6362_n6133) );
	NAND2X1 NAND2X1_4259 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6131), .B(dp.rf._abc_6362_n6133), .Y(dp.rf._abc_6362_n6134) );
	NAND2X1 NAND2X1_4260 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<7>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6135) );
	NAND2X1 NAND2X1_4261 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<7>), .Y(dp.rf._abc_6362_n6136) );
	AND2X2 AND2X2_138 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6136), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6137) );
	NAND2X1 NAND2X1_4262 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6135), .B(dp.rf._abc_6362_n6137), .Y(dp.rf._abc_6362_n6138) );
	NAND2X1 NAND2X1_4263 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6134), .B(dp.rf._abc_6362_n6138), .Y(dp.rf._abc_6362_n6139) );
	AND2X2 AND2X2_139 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6139), .B(instr[23]), .Y(dp.rf._abc_6362_n6140) );
	NAND2X1 NAND2X1_4264 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<7>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6141) );
	NAND2X1 NAND2X1_4265 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<7>), .Y(dp.rf._abc_6362_n6142) );
	AND2X2 AND2X2_140 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6142), .B(instr[22]), .Y(dp.rf._abc_6362_n6143) );
	NAND2X1 NAND2X1_4266 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6141), .B(dp.rf._abc_6362_n6143), .Y(dp.rf._abc_6362_n6144) );
	NAND2X1 NAND2X1_4267 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<7>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6145) );
	NAND2X1 NAND2X1_4268 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<7>), .Y(dp.rf._abc_6362_n6146) );
	AND2X2 AND2X2_141 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6146), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6147) );
	NAND2X1 NAND2X1_4269 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6145), .B(dp.rf._abc_6362_n6147), .Y(dp.rf._abc_6362_n6148) );
	NAND2X1 NAND2X1_4270 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6144), .B(dp.rf._abc_6362_n6148), .Y(dp.rf._abc_6362_n6149) );
	NAND2X1 NAND2X1_4271 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6149), .Y(dp.rf._abc_6362_n6150) );
	NAND2X1 NAND2X1_4272 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6150), .Y(dp.rf._abc_6362_n6151) );
	NOR2X1 NOR2X1_402 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6140), .B(dp.rf._abc_6362_n6151), .Y(dp.rf._abc_6362_n6152) );
	NOR2X1 NOR2X1_403 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6152), .Y(dp.rf._abc_6362_n6153) );
	NAND2X1 NAND2X1_4273 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6130), .B(dp.rf._abc_6362_n6153), .Y(dp.rf._abc_6362_n6154) );
	NAND2X1 NAND2X1_4274 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n6154), .Y(dp.rf._abc_6362_n6155) );
	NOR2X1 NOR2X1_404 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6104), .B(dp.rf._abc_6362_n6155), .Y(dp.srca_7_) );
	NAND2X1 NAND2X1_4275 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<8>), .Y(dp.rf._abc_6362_n6157) );
	NAND2X1 NAND2X1_4276 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6158) );
	NAND2X1 NAND2X1_4277 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6157), .B(dp.rf._abc_6362_n6158), .Y(dp.rf._abc_6362_n6159) );
	NAND2X1 NAND2X1_4278 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6159), .Y(dp.rf._abc_6362_n6160) );
	NAND2X1 NAND2X1_4279 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<8>), .Y(dp.rf._abc_6362_n6161) );
	NAND2X1 NAND2X1_4280 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6162) );
	NAND2X1 NAND2X1_4281 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6161), .B(dp.rf._abc_6362_n6162), .Y(dp.rf._abc_6362_n6163) );
	NAND2X1 NAND2X1_4282 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6163), .Y(dp.rf._abc_6362_n6164) );
	NAND2X1 NAND2X1_4283 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6160), .B(dp.rf._abc_6362_n6164), .Y(dp.rf._abc_6362_n6165) );
	NOR2X1 NOR2X1_405 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6165), .Y(dp.rf._abc_6362_n6166) );
	NAND2X1 NAND2X1_4284 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<8>), .Y(dp.rf._abc_6362_n6167) );
	NAND2X1 NAND2X1_4285 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6168) );
	NAND2X1 NAND2X1_4286 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6167), .B(dp.rf._abc_6362_n6168), .Y(dp.rf._abc_6362_n6169) );
	NAND2X1 NAND2X1_4287 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6169), .Y(dp.rf._abc_6362_n6170) );
	NAND2X1 NAND2X1_4288 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<8>), .Y(dp.rf._abc_6362_n6171) );
	NAND2X1 NAND2X1_4289 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6172) );
	NAND2X1 NAND2X1_4290 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6171), .B(dp.rf._abc_6362_n6172), .Y(dp.rf._abc_6362_n6173) );
	NAND2X1 NAND2X1_4291 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6173), .Y(dp.rf._abc_6362_n6174) );
	AND2X2 AND2X2_142 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6170), .B(dp.rf._abc_6362_n6174), .Y(dp.rf._abc_6362_n6175) );
	NAND2X1 NAND2X1_4292 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6175), .Y(dp.rf._abc_6362_n6176) );
	NAND2X1 NAND2X1_4293 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n6176), .Y(dp.rf._abc_6362_n6177) );
	NOR2X1 NOR2X1_406 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6166), .B(dp.rf._abc_6362_n6177), .Y(dp.rf._abc_6362_n6178) );
	NAND2X1 NAND2X1_4294 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<8>), .Y(dp.rf._abc_6362_n6179) );
	NAND2X1 NAND2X1_4295 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6179), .Y(dp.rf._abc_6362_n6180) );
	INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<8>), .Y(dp.rf._abc_6362_n6181) );
	NOR2X1 NOR2X1_407 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6181), .Y(dp.rf._abc_6362_n6182) );
	NOR2X1 NOR2X1_408 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6180), .B(dp.rf._abc_6362_n6182), .Y(dp.rf._abc_6362_n6183) );
	NAND2X1 NAND2X1_4296 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<8>), .Y(dp.rf._abc_6362_n6184) );
	NAND2X1 NAND2X1_4297 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6184), .Y(dp.rf._abc_6362_n6185) );
	INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<8>), .Y(dp.rf._abc_6362_n6186) );
	NOR2X1 NOR2X1_409 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6186), .Y(dp.rf._abc_6362_n6187) );
	NOR2X1 NOR2X1_410 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6185), .B(dp.rf._abc_6362_n6187), .Y(dp.rf._abc_6362_n6188) );
	NOR2X1 NOR2X1_411 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6183), .B(dp.rf._abc_6362_n6188), .Y(dp.rf._abc_6362_n6189) );
	NAND2X1 NAND2X1_4298 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6189), .Y(dp.rf._abc_6362_n6190) );
	NAND2X1 NAND2X1_4299 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<8>), .Y(dp.rf._abc_6362_n6191) );
	NAND2X1 NAND2X1_4300 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6191), .Y(dp.rf._abc_6362_n6192) );
	INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<8>), .Y(dp.rf._abc_6362_n6193) );
	NOR2X1 NOR2X1_412 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6193), .Y(dp.rf._abc_6362_n6194) );
	NOR2X1 NOR2X1_413 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6192), .B(dp.rf._abc_6362_n6194), .Y(dp.rf._abc_6362_n6195) );
	NAND2X1 NAND2X1_4301 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<8>), .Y(dp.rf._abc_6362_n6196) );
	NAND2X1 NAND2X1_4302 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6196), .Y(dp.rf._abc_6362_n6197) );
	INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<8>), .Y(dp.rf._abc_6362_n6198) );
	NOR2X1 NOR2X1_414 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6198), .Y(dp.rf._abc_6362_n6199) );
	NOR2X1 NOR2X1_415 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6197), .B(dp.rf._abc_6362_n6199), .Y(dp.rf._abc_6362_n6200) );
	NOR2X1 NOR2X1_416 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6195), .B(dp.rf._abc_6362_n6200), .Y(dp.rf._abc_6362_n6201) );
	NAND2X1 NAND2X1_4303 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6201), .Y(dp.rf._abc_6362_n6202) );
	NAND2X1 NAND2X1_4304 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6190), .B(dp.rf._abc_6362_n6202), .Y(dp.rf._abc_6362_n6203) );
	NAND2X1 NAND2X1_4305 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6203), .Y(dp.rf._abc_6362_n6204) );
	NAND2X1 NAND2X1_4306 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6204), .Y(dp.rf._abc_6362_n6205) );
	NOR2X1 NOR2X1_417 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6178), .B(dp.rf._abc_6362_n6205), .Y(dp.rf._abc_6362_n6206) );
	NAND2X1 NAND2X1_4307 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<8>), .Y(dp.rf._abc_6362_n6207) );
	NAND2X1 NAND2X1_4308 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6208) );
	NAND2X1 NAND2X1_4309 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6207), .B(dp.rf._abc_6362_n6208), .Y(dp.rf._abc_6362_n6209) );
	NAND2X1 NAND2X1_4310 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6209), .Y(dp.rf._abc_6362_n6210) );
	NAND2X1 NAND2X1_4311 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<8>), .Y(dp.rf._abc_6362_n6211) );
	NAND2X1 NAND2X1_4312 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6212) );
	NAND2X1 NAND2X1_4313 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6211), .B(dp.rf._abc_6362_n6212), .Y(dp.rf._abc_6362_n6213) );
	NAND2X1 NAND2X1_4314 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6213), .Y(dp.rf._abc_6362_n6214) );
	AND2X2 AND2X2_143 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6210), .B(dp.rf._abc_6362_n6214), .Y(dp.rf._abc_6362_n6215) );
	NAND2X1 NAND2X1_4315 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6215), .Y(dp.rf._abc_6362_n6216) );
	NAND2X1 NAND2X1_4316 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<8>), .Y(dp.rf._abc_6362_n6217) );
	NAND2X1 NAND2X1_4317 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6218) );
	NAND2X1 NAND2X1_4318 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6217), .B(dp.rf._abc_6362_n6218), .Y(dp.rf._abc_6362_n6219) );
	NAND2X1 NAND2X1_4319 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6219), .Y(dp.rf._abc_6362_n6220) );
	NAND2X1 NAND2X1_4320 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<8>), .Y(dp.rf._abc_6362_n6221) );
	NAND2X1 NAND2X1_4321 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6222) );
	NAND2X1 NAND2X1_4322 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6221), .B(dp.rf._abc_6362_n6222), .Y(dp.rf._abc_6362_n6223) );
	NAND2X1 NAND2X1_4323 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6223), .Y(dp.rf._abc_6362_n6224) );
	AND2X2 AND2X2_144 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6220), .B(dp.rf._abc_6362_n6224), .Y(dp.rf._abc_6362_n6225) );
	NAND2X1 NAND2X1_4324 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6225), .Y(dp.rf._abc_6362_n6226) );
	AND2X2 AND2X2_145 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6226), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n6227) );
	NAND2X1 NAND2X1_4325 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6216), .B(dp.rf._abc_6362_n6227), .Y(dp.rf._abc_6362_n6228) );
	NAND2X1 NAND2X1_4326 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6229) );
	NAND2X1 NAND2X1_4327 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<8>), .Y(dp.rf._abc_6362_n6230) );
	AND2X2 AND2X2_146 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6230), .B(instr[22]), .Y(dp.rf._abc_6362_n6231) );
	NAND2X1 NAND2X1_4328 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6229), .B(dp.rf._abc_6362_n6231), .Y(dp.rf._abc_6362_n6232) );
	NAND2X1 NAND2X1_4329 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6233) );
	NAND2X1 NAND2X1_4330 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<8>), .Y(dp.rf._abc_6362_n6234) );
	AND2X2 AND2X2_147 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6234), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6235) );
	NAND2X1 NAND2X1_4331 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6233), .B(dp.rf._abc_6362_n6235), .Y(dp.rf._abc_6362_n6236) );
	NAND2X1 NAND2X1_4332 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6232), .B(dp.rf._abc_6362_n6236), .Y(dp.rf._abc_6362_n6237) );
	AND2X2 AND2X2_148 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6237), .B(instr[23]), .Y(dp.rf._abc_6362_n6238) );
	NAND2X1 NAND2X1_4333 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6239) );
	NAND2X1 NAND2X1_4334 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<8>), .Y(dp.rf._abc_6362_n6240) );
	AND2X2 AND2X2_149 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6240), .B(instr[22]), .Y(dp.rf._abc_6362_n6241) );
	NAND2X1 NAND2X1_4335 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6239), .B(dp.rf._abc_6362_n6241), .Y(dp.rf._abc_6362_n6242) );
	NAND2X1 NAND2X1_4336 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<8>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6243) );
	NAND2X1 NAND2X1_4337 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<8>), .Y(dp.rf._abc_6362_n6244) );
	AND2X2 AND2X2_150 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6244), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6245) );
	NAND2X1 NAND2X1_4338 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6243), .B(dp.rf._abc_6362_n6245), .Y(dp.rf._abc_6362_n6246) );
	NAND2X1 NAND2X1_4339 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6242), .B(dp.rf._abc_6362_n6246), .Y(dp.rf._abc_6362_n6247) );
	NAND2X1 NAND2X1_4340 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6247), .Y(dp.rf._abc_6362_n6248) );
	NAND2X1 NAND2X1_4341 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6248), .Y(dp.rf._abc_6362_n6249) );
	NOR2X1 NOR2X1_418 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6238), .B(dp.rf._abc_6362_n6249), .Y(dp.rf._abc_6362_n6250) );
	NOR2X1 NOR2X1_419 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6250), .Y(dp.rf._abc_6362_n6251) );
	NAND2X1 NAND2X1_4342 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6228), .B(dp.rf._abc_6362_n6251), .Y(dp.rf._abc_6362_n6252) );
	NAND2X1 NAND2X1_4343 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n6252), .Y(dp.rf._abc_6362_n6253) );
	NOR2X1 NOR2X1_420 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6206), .B(dp.rf._abc_6362_n6253), .Y(dp.srca_8_) );
	NAND2X1 NAND2X1_4344 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<9>), .Y(dp.rf._abc_6362_n6255) );
	NAND2X1 NAND2X1_4345 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6255), .Y(dp.rf._abc_6362_n6256) );
	INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<9>), .Y(dp.rf._abc_6362_n6257) );
	NOR2X1 NOR2X1_421 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6257), .Y(dp.rf._abc_6362_n6258) );
	NOR2X1 NOR2X1_422 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6256), .B(dp.rf._abc_6362_n6258), .Y(dp.rf._abc_6362_n6259) );
	NAND2X1 NAND2X1_4346 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<9>), .Y(dp.rf._abc_6362_n6260) );
	NAND2X1 NAND2X1_4347 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6260), .Y(dp.rf._abc_6362_n6261) );
	INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<9>), .Y(dp.rf._abc_6362_n6262) );
	NOR2X1 NOR2X1_423 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6262), .Y(dp.rf._abc_6362_n6263) );
	NOR2X1 NOR2X1_424 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6261), .B(dp.rf._abc_6362_n6263), .Y(dp.rf._abc_6362_n6264) );
	NOR2X1 NOR2X1_425 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6259), .B(dp.rf._abc_6362_n6264), .Y(dp.rf._abc_6362_n6265) );
	NAND2X1 NAND2X1_4348 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6265), .Y(dp.rf._abc_6362_n6266) );
	NAND2X1 NAND2X1_4349 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<9>), .Y(dp.rf._abc_6362_n6267) );
	NAND2X1 NAND2X1_4350 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6267), .Y(dp.rf._abc_6362_n6268) );
	INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<9>), .Y(dp.rf._abc_6362_n6269) );
	NOR2X1 NOR2X1_426 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6269), .Y(dp.rf._abc_6362_n6270) );
	NOR2X1 NOR2X1_427 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6268), .B(dp.rf._abc_6362_n6270), .Y(dp.rf._abc_6362_n6271) );
	NAND2X1 NAND2X1_4351 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<9>), .Y(dp.rf._abc_6362_n6272) );
	NAND2X1 NAND2X1_4352 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6272), .Y(dp.rf._abc_6362_n6273) );
	INVX1 INVX1_113 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<9>), .Y(dp.rf._abc_6362_n6274) );
	NOR2X1 NOR2X1_428 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6274), .Y(dp.rf._abc_6362_n6275) );
	NOR2X1 NOR2X1_429 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6273), .B(dp.rf._abc_6362_n6275), .Y(dp.rf._abc_6362_n6276) );
	NOR2X1 NOR2X1_430 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6271), .B(dp.rf._abc_6362_n6276), .Y(dp.rf._abc_6362_n6277) );
	NAND2X1 NAND2X1_4353 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6277), .Y(dp.rf._abc_6362_n6278) );
	NAND2X1 NAND2X1_4354 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6266), .B(dp.rf._abc_6362_n6278), .Y(dp.rf._abc_6362_n6279) );
	NAND2X1 NAND2X1_4355 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6279), .Y(dp.rf._abc_6362_n6280) );
	NAND2X1 NAND2X1_4356 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<9>), .Y(dp.rf._abc_6362_n6281) );
	NAND2X1 NAND2X1_4357 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6281), .Y(dp.rf._abc_6362_n6282) );
	INVX1 INVX1_114 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<9>), .Y(dp.rf._abc_6362_n6283) );
	NOR2X1 NOR2X1_431 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6283), .Y(dp.rf._abc_6362_n6284) );
	NOR2X1 NOR2X1_432 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6282), .B(dp.rf._abc_6362_n6284), .Y(dp.rf._abc_6362_n6285) );
	NAND2X1 NAND2X1_4358 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<9>), .Y(dp.rf._abc_6362_n6286) );
	NAND2X1 NAND2X1_4359 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6286), .Y(dp.rf._abc_6362_n6287) );
	INVX1 INVX1_115 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<9>), .Y(dp.rf._abc_6362_n6288) );
	NOR2X1 NOR2X1_433 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6288), .Y(dp.rf._abc_6362_n6289) );
	NOR2X1 NOR2X1_434 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6287), .B(dp.rf._abc_6362_n6289), .Y(dp.rf._abc_6362_n6290) );
	OR2X2 OR2X2_42 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6285), .B(dp.rf._abc_6362_n6290), .Y(dp.rf._abc_6362_n6291) );
	NAND2X1 NAND2X1_4360 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6291), .Y(dp.rf._abc_6362_n6292) );
	NAND2X1 NAND2X1_4361 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<9>), .Y(dp.rf._abc_6362_n6293) );
	NAND2X1 NAND2X1_4362 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6293), .Y(dp.rf._abc_6362_n6294) );
	INVX1 INVX1_116 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<9>), .Y(dp.rf._abc_6362_n6295) );
	NOR2X1 NOR2X1_435 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6295), .Y(dp.rf._abc_6362_n6296) );
	NOR2X1 NOR2X1_436 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6294), .B(dp.rf._abc_6362_n6296), .Y(dp.rf._abc_6362_n6297) );
	NAND2X1 NAND2X1_4363 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<9>), .Y(dp.rf._abc_6362_n6298) );
	NAND2X1 NAND2X1_4364 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6298), .Y(dp.rf._abc_6362_n6299) );
	INVX1 INVX1_117 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<9>), .Y(dp.rf._abc_6362_n6300) );
	NOR2X1 NOR2X1_437 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6300), .Y(dp.rf._abc_6362_n6301) );
	NOR2X1 NOR2X1_438 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6299), .B(dp.rf._abc_6362_n6301), .Y(dp.rf._abc_6362_n6302) );
	OR2X2 OR2X2_43 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6297), .B(dp.rf._abc_6362_n6302), .Y(dp.rf._abc_6362_n6303) );
	NAND2X1 NAND2X1_4365 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6303), .Y(dp.rf._abc_6362_n6304) );
	AND2X2 AND2X2_151 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6304), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n6305) );
	NAND2X1 NAND2X1_4366 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6292), .B(dp.rf._abc_6362_n6305), .Y(dp.rf._abc_6362_n6306) );
	NAND2X1 NAND2X1_4367 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6280), .B(dp.rf._abc_6362_n6306), .Y(dp.rf._abc_6362_n6307) );
	NOR2X1 NOR2X1_439 ( .gnd(gnd), .vdd(vdd), .A(instr[25]), .B(dp.rf._abc_6362_n6307), .Y(dp.rf._abc_6362_n6308) );
	NAND2X1 NAND2X1_4368 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<9>), .Y(dp.rf._abc_6362_n6309) );
	NAND2X1 NAND2X1_4369 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<9>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6310) );
	NAND2X1 NAND2X1_4370 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6309), .B(dp.rf._abc_6362_n6310), .Y(dp.rf._abc_6362_n6311) );
	NAND2X1 NAND2X1_4371 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6311), .Y(dp.rf._abc_6362_n6312) );
	NAND2X1 NAND2X1_4372 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<9>), .Y(dp.rf._abc_6362_n6313) );
	NAND2X1 NAND2X1_4373 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<9>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6314) );
	NAND2X1 NAND2X1_4374 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6313), .B(dp.rf._abc_6362_n6314), .Y(dp.rf._abc_6362_n6315) );
	NAND2X1 NAND2X1_4375 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6315), .Y(dp.rf._abc_6362_n6316) );
	AND2X2 AND2X2_152 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6312), .B(dp.rf._abc_6362_n6316), .Y(dp.rf._abc_6362_n6317) );
	NAND2X1 NAND2X1_4376 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6317), .Y(dp.rf._abc_6362_n6318) );
	NAND2X1 NAND2X1_4377 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<9>), .Y(dp.rf._abc_6362_n6319) );
	NAND2X1 NAND2X1_4378 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<9>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6320) );
	NAND2X1 NAND2X1_4379 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6319), .B(dp.rf._abc_6362_n6320), .Y(dp.rf._abc_6362_n6321) );
	NAND2X1 NAND2X1_4380 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6321), .Y(dp.rf._abc_6362_n6322) );
	NAND2X1 NAND2X1_4381 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<9>), .Y(dp.rf._abc_6362_n6323) );
	NAND2X1 NAND2X1_4382 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<9>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6324) );
	NAND2X1 NAND2X1_4383 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6323), .B(dp.rf._abc_6362_n6324), .Y(dp.rf._abc_6362_n6325) );
	NAND2X1 NAND2X1_4384 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6325), .Y(dp.rf._abc_6362_n6326) );
	AND2X2 AND2X2_153 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6322), .B(dp.rf._abc_6362_n6326), .Y(dp.rf._abc_6362_n6327) );
	NAND2X1 NAND2X1_4385 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6327), .Y(dp.rf._abc_6362_n6328) );
	AND2X2 AND2X2_154 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6328), .B(instr[24]), .Y(dp.rf._abc_6362_n6329) );
	NAND2X1 NAND2X1_4386 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6318), .B(dp.rf._abc_6362_n6329), .Y(dp.rf._abc_6362_n6330) );
	NAND2X1 NAND2X1_4387 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<9>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6331) );
	NAND2X1 NAND2X1_4388 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<9>), .Y(dp.rf._abc_6362_n6332) );
	AND2X2 AND2X2_155 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6332), .B(instr[22]), .Y(dp.rf._abc_6362_n6333) );
	NAND2X1 NAND2X1_4389 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6331), .B(dp.rf._abc_6362_n6333), .Y(dp.rf._abc_6362_n6334) );
	NAND2X1 NAND2X1_4390 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<9>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6335) );
	NAND2X1 NAND2X1_4391 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<9>), .Y(dp.rf._abc_6362_n6336) );
	AND2X2 AND2X2_156 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6336), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6337) );
	NAND2X1 NAND2X1_4392 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6335), .B(dp.rf._abc_6362_n6337), .Y(dp.rf._abc_6362_n6338) );
	NAND2X1 NAND2X1_4393 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6334), .B(dp.rf._abc_6362_n6338), .Y(dp.rf._abc_6362_n6339) );
	AND2X2 AND2X2_157 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6339), .B(instr[23]), .Y(dp.rf._abc_6362_n6340) );
	NAND2X1 NAND2X1_4394 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<9>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6341) );
	NAND2X1 NAND2X1_4395 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<9>), .Y(dp.rf._abc_6362_n6342) );
	AND2X2 AND2X2_158 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6342), .B(instr[22]), .Y(dp.rf._abc_6362_n6343) );
	NAND2X1 NAND2X1_4396 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6341), .B(dp.rf._abc_6362_n6343), .Y(dp.rf._abc_6362_n6344) );
	NAND2X1 NAND2X1_4397 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<9>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6345) );
	NAND2X1 NAND2X1_4398 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<9>), .Y(dp.rf._abc_6362_n6346) );
	AND2X2 AND2X2_159 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6346), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6347) );
	NAND2X1 NAND2X1_4399 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6345), .B(dp.rf._abc_6362_n6347), .Y(dp.rf._abc_6362_n6348) );
	NAND2X1 NAND2X1_4400 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6344), .B(dp.rf._abc_6362_n6348), .Y(dp.rf._abc_6362_n6349) );
	NAND2X1 NAND2X1_4401 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6349), .Y(dp.rf._abc_6362_n6350) );
	NAND2X1 NAND2X1_4402 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n6350), .Y(dp.rf._abc_6362_n6351) );
	NOR2X1 NOR2X1_440 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6340), .B(dp.rf._abc_6362_n6351), .Y(dp.rf._abc_6362_n6352) );
	NOR2X1 NOR2X1_441 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6352), .Y(dp.rf._abc_6362_n6353) );
	NAND2X1 NAND2X1_4403 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6330), .B(dp.rf._abc_6362_n6353), .Y(dp.rf._abc_6362_n6354) );
	NAND2X1 NAND2X1_4404 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n6354), .Y(dp.rf._abc_6362_n6355) );
	NOR2X1 NOR2X1_442 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6308), .B(dp.rf._abc_6362_n6355), .Y(dp.srca_9_) );
	NAND2X1 NAND2X1_4405 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<10>), .Y(dp.rf._abc_6362_n6357) );
	NAND2X1 NAND2X1_4406 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6357), .Y(dp.rf._abc_6362_n6358) );
	INVX1 INVX1_118 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<10>), .Y(dp.rf._abc_6362_n6359) );
	NOR2X1 NOR2X1_443 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6359), .Y(dp.rf._abc_6362_n6360) );
	NOR2X1 NOR2X1_444 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6358), .B(dp.rf._abc_6362_n6360), .Y(dp.rf._abc_6362_n6361) );
	NAND2X1 NAND2X1_4407 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<10>), .Y(dp.rf._abc_6362_n6362) );
	NAND2X1 NAND2X1_4408 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6362), .Y(dp.rf._abc_6362_n6363) );
	INVX1 INVX1_119 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<10>), .Y(dp.rf._abc_6362_n6364) );
	NOR2X1 NOR2X1_445 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6364), .Y(dp.rf._abc_6362_n6365) );
	NOR2X1 NOR2X1_446 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6363), .B(dp.rf._abc_6362_n6365), .Y(dp.rf._abc_6362_n6366) );
	NOR2X1 NOR2X1_447 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6361), .B(dp.rf._abc_6362_n6366), .Y(dp.rf._abc_6362_n6367) );
	NAND2X1 NAND2X1_4409 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6367), .Y(dp.rf._abc_6362_n6368) );
	NAND2X1 NAND2X1_4410 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<10>), .Y(dp.rf._abc_6362_n6369) );
	NAND2X1 NAND2X1_4411 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6369), .Y(dp.rf._abc_6362_n6370) );
	INVX1 INVX1_120 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<10>), .Y(dp.rf._abc_6362_n6371) );
	NOR2X1 NOR2X1_448 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6371), .Y(dp.rf._abc_6362_n6372) );
	NOR2X1 NOR2X1_449 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6370), .B(dp.rf._abc_6362_n6372), .Y(dp.rf._abc_6362_n6373) );
	NAND2X1 NAND2X1_4412 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<10>), .Y(dp.rf._abc_6362_n6374) );
	NAND2X1 NAND2X1_4413 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6374), .Y(dp.rf._abc_6362_n6375) );
	INVX1 INVX1_121 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<10>), .Y(dp.rf._abc_6362_n6376) );
	NOR2X1 NOR2X1_450 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6376), .Y(dp.rf._abc_6362_n6377) );
	NOR2X1 NOR2X1_451 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6375), .B(dp.rf._abc_6362_n6377), .Y(dp.rf._abc_6362_n6378) );
	NOR2X1 NOR2X1_452 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6373), .B(dp.rf._abc_6362_n6378), .Y(dp.rf._abc_6362_n6379) );
	NAND2X1 NAND2X1_4414 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6379), .Y(dp.rf._abc_6362_n6380) );
	NAND2X1 NAND2X1_4415 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6368), .B(dp.rf._abc_6362_n6380), .Y(dp.rf._abc_6362_n6381) );
	NAND2X1 NAND2X1_4416 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6381), .Y(dp.rf._abc_6362_n6382) );
	NAND2X1 NAND2X1_4417 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<10>), .Y(dp.rf._abc_6362_n6383) );
	NAND2X1 NAND2X1_4418 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<10>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6384) );
	NAND2X1 NAND2X1_4419 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6383), .B(dp.rf._abc_6362_n6384), .Y(dp.rf._abc_6362_n6385) );
	NAND2X1 NAND2X1_4420 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6385), .Y(dp.rf._abc_6362_n6386) );
	NAND2X1 NAND2X1_4421 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<10>), .Y(dp.rf._abc_6362_n6387) );
	NAND2X1 NAND2X1_4422 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<10>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6388) );
	NAND2X1 NAND2X1_4423 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6387), .B(dp.rf._abc_6362_n6388), .Y(dp.rf._abc_6362_n6389) );
	NAND2X1 NAND2X1_4424 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6389), .Y(dp.rf._abc_6362_n6390) );
	AND2X2 AND2X2_160 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6386), .B(dp.rf._abc_6362_n6390), .Y(dp.rf._abc_6362_n6391) );
	NAND2X1 NAND2X1_4425 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6391), .Y(dp.rf._abc_6362_n6392) );
	NAND2X1 NAND2X1_4426 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<10>), .Y(dp.rf._abc_6362_n6393) );
	NAND2X1 NAND2X1_4427 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6393), .Y(dp.rf._abc_6362_n6394) );
	AND2X2 AND2X2_161 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf.rf_2_<10>), .Y(dp.rf._abc_6362_n6395) );
	NOR2X1 NOR2X1_453 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6394), .B(dp.rf._abc_6362_n6395), .Y(dp.rf._abc_6362_n6396) );
	NAND2X1 NAND2X1_4428 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<10>), .Y(dp.rf._abc_6362_n6397) );
	NAND2X1 NAND2X1_4429 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6397), .Y(dp.rf._abc_6362_n6398) );
	INVX1 INVX1_122 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<10>), .Y(dp.rf._abc_6362_n6399) );
	NOR2X1 NOR2X1_454 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6399), .Y(dp.rf._abc_6362_n6400) );
	NOR2X1 NOR2X1_455 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6398), .B(dp.rf._abc_6362_n6400), .Y(dp.rf._abc_6362_n6401) );
	OR2X2 OR2X2_44 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6396), .B(dp.rf._abc_6362_n6401), .Y(dp.rf._abc_6362_n6402) );
	NAND2X1 NAND2X1_4430 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6402), .Y(dp.rf._abc_6362_n6403) );
	AND2X2 AND2X2_162 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6403), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n6404) );
	NAND2X1 NAND2X1_4431 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6392), .B(dp.rf._abc_6362_n6404), .Y(dp.rf._abc_6362_n6405) );
	NAND2X1 NAND2X1_4432 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6382), .B(dp.rf._abc_6362_n6405), .Y(dp.rf._abc_6362_n6406) );
	NOR2X1 NOR2X1_456 ( .gnd(gnd), .vdd(vdd), .A(instr[25]), .B(dp.rf._abc_6362_n6406), .Y(dp.rf._abc_6362_n6407) );
	NAND2X1 NAND2X1_4433 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<10>), .Y(dp.rf._abc_6362_n6408) );
	NAND2X1 NAND2X1_4434 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6408), .Y(dp.rf._abc_6362_n6409) );
	INVX1 INVX1_123 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<10>), .Y(dp.rf._abc_6362_n6410) );
	NOR2X1 NOR2X1_457 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6410), .Y(dp.rf._abc_6362_n6411) );
	NOR2X1 NOR2X1_458 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6409), .B(dp.rf._abc_6362_n6411), .Y(dp.rf._abc_6362_n6412) );
	NAND2X1 NAND2X1_4435 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<10>), .Y(dp.rf._abc_6362_n6413) );
	NAND2X1 NAND2X1_4436 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6413), .Y(dp.rf._abc_6362_n6414) );
	INVX1 INVX1_124 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<10>), .Y(dp.rf._abc_6362_n6415) );
	NOR2X1 NOR2X1_459 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6415), .Y(dp.rf._abc_6362_n6416) );
	NOR2X1 NOR2X1_460 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6414), .B(dp.rf._abc_6362_n6416), .Y(dp.rf._abc_6362_n6417) );
	OR2X2 OR2X2_45 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6412), .B(dp.rf._abc_6362_n6417), .Y(dp.rf._abc_6362_n6418) );
	NAND2X1 NAND2X1_4437 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6418), .Y(dp.rf._abc_6362_n6419) );
	NAND2X1 NAND2X1_4438 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<10>), .Y(dp.rf._abc_6362_n6420) );
	NAND2X1 NAND2X1_4439 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6420), .Y(dp.rf._abc_6362_n6421) );
	INVX1 INVX1_125 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<10>), .Y(dp.rf._abc_6362_n6422) );
	NOR2X1 NOR2X1_461 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6422), .Y(dp.rf._abc_6362_n6423) );
	NOR2X1 NOR2X1_462 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6421), .B(dp.rf._abc_6362_n6423), .Y(dp.rf._abc_6362_n6424) );
	NAND2X1 NAND2X1_4440 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<10>), .Y(dp.rf._abc_6362_n6425) );
	NAND2X1 NAND2X1_4441 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6425), .Y(dp.rf._abc_6362_n6426) );
	INVX1 INVX1_126 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<10>), .Y(dp.rf._abc_6362_n6427) );
	NOR2X1 NOR2X1_463 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6427), .Y(dp.rf._abc_6362_n6428) );
	NOR2X1 NOR2X1_464 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6426), .B(dp.rf._abc_6362_n6428), .Y(dp.rf._abc_6362_n6429) );
	OR2X2 OR2X2_46 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6424), .B(dp.rf._abc_6362_n6429), .Y(dp.rf._abc_6362_n6430) );
	NAND2X1 NAND2X1_4442 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6430), .Y(dp.rf._abc_6362_n6431) );
	AND2X2 AND2X2_163 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6431), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n6432) );
	NAND2X1 NAND2X1_4443 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6419), .B(dp.rf._abc_6362_n6432), .Y(dp.rf._abc_6362_n6433) );
	NAND2X1 NAND2X1_4444 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<10>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6434) );
	NAND2X1 NAND2X1_4445 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<10>), .Y(dp.rf._abc_6362_n6435) );
	AND2X2 AND2X2_164 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6435), .B(instr[22]), .Y(dp.rf._abc_6362_n6436) );
	NAND2X1 NAND2X1_4446 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6434), .B(dp.rf._abc_6362_n6436), .Y(dp.rf._abc_6362_n6437) );
	NAND2X1 NAND2X1_4447 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<10>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6438) );
	NAND2X1 NAND2X1_4448 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<10>), .Y(dp.rf._abc_6362_n6439) );
	AND2X2 AND2X2_165 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6439), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6440) );
	NAND2X1 NAND2X1_4449 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6438), .B(dp.rf._abc_6362_n6440), .Y(dp.rf._abc_6362_n6441) );
	NAND2X1 NAND2X1_4450 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6437), .B(dp.rf._abc_6362_n6441), .Y(dp.rf._abc_6362_n6442) );
	AND2X2 AND2X2_166 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6442), .B(instr[23]), .Y(dp.rf._abc_6362_n6443) );
	NAND2X1 NAND2X1_4451 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<10>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6444) );
	NAND2X1 NAND2X1_4452 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<10>), .Y(dp.rf._abc_6362_n6445) );
	AND2X2 AND2X2_167 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6445), .B(instr[22]), .Y(dp.rf._abc_6362_n6446) );
	NAND2X1 NAND2X1_4453 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6444), .B(dp.rf._abc_6362_n6446), .Y(dp.rf._abc_6362_n6447) );
	NAND2X1 NAND2X1_4454 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<10>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6448) );
	NAND2X1 NAND2X1_4455 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<10>), .Y(dp.rf._abc_6362_n6449) );
	AND2X2 AND2X2_168 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6449), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6450) );
	NAND2X1 NAND2X1_4456 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6448), .B(dp.rf._abc_6362_n6450), .Y(dp.rf._abc_6362_n6451) );
	NAND2X1 NAND2X1_4457 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6447), .B(dp.rf._abc_6362_n6451), .Y(dp.rf._abc_6362_n6452) );
	NAND2X1 NAND2X1_4458 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6452), .Y(dp.rf._abc_6362_n6453) );
	NAND2X1 NAND2X1_4459 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6453), .Y(dp.rf._abc_6362_n6454) );
	NOR2X1 NOR2X1_465 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6443), .B(dp.rf._abc_6362_n6454), .Y(dp.rf._abc_6362_n6455) );
	NOR2X1 NOR2X1_466 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6455), .Y(dp.rf._abc_6362_n6456) );
	NAND2X1 NAND2X1_4460 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6433), .B(dp.rf._abc_6362_n6456), .Y(dp.rf._abc_6362_n6457) );
	NAND2X1 NAND2X1_4461 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n6457), .Y(dp.rf._abc_6362_n6458) );
	NOR2X1 NOR2X1_467 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6407), .B(dp.rf._abc_6362_n6458), .Y(dp.srca_10_) );
	NAND2X1 NAND2X1_4462 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<11>), .Y(dp.rf._abc_6362_n6460) );
	NAND2X1 NAND2X1_4463 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6460), .Y(dp.rf._abc_6362_n6461) );
	INVX1 INVX1_127 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<11>), .Y(dp.rf._abc_6362_n6462) );
	NOR2X1 NOR2X1_468 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6462), .Y(dp.rf._abc_6362_n6463) );
	NOR2X1 NOR2X1_469 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6461), .B(dp.rf._abc_6362_n6463), .Y(dp.rf._abc_6362_n6464) );
	NAND2X1 NAND2X1_4464 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<11>), .Y(dp.rf._abc_6362_n6465) );
	NAND2X1 NAND2X1_4465 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6465), .Y(dp.rf._abc_6362_n6466) );
	INVX1 INVX1_128 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<11>), .Y(dp.rf._abc_6362_n6467) );
	NOR2X1 NOR2X1_470 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6467), .Y(dp.rf._abc_6362_n6468) );
	NOR2X1 NOR2X1_471 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6466), .B(dp.rf._abc_6362_n6468), .Y(dp.rf._abc_6362_n6469) );
	NOR2X1 NOR2X1_472 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6464), .B(dp.rf._abc_6362_n6469), .Y(dp.rf._abc_6362_n6470) );
	NAND2X1 NAND2X1_4466 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6470), .Y(dp.rf._abc_6362_n6471) );
	NAND2X1 NAND2X1_4467 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<11>), .Y(dp.rf._abc_6362_n6472) );
	NAND2X1 NAND2X1_4468 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6472), .Y(dp.rf._abc_6362_n6473) );
	INVX1 INVX1_129 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<11>), .Y(dp.rf._abc_6362_n6474) );
	NOR2X1 NOR2X1_473 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6474), .Y(dp.rf._abc_6362_n6475) );
	NOR2X1 NOR2X1_474 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6473), .B(dp.rf._abc_6362_n6475), .Y(dp.rf._abc_6362_n6476) );
	NAND2X1 NAND2X1_4469 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<11>), .Y(dp.rf._abc_6362_n6477) );
	NAND2X1 NAND2X1_4470 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6477), .Y(dp.rf._abc_6362_n6478) );
	INVX1 INVX1_130 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<11>), .Y(dp.rf._abc_6362_n6479) );
	NOR2X1 NOR2X1_475 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6479), .Y(dp.rf._abc_6362_n6480) );
	NOR2X1 NOR2X1_476 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6478), .B(dp.rf._abc_6362_n6480), .Y(dp.rf._abc_6362_n6481) );
	NOR2X1 NOR2X1_477 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6476), .B(dp.rf._abc_6362_n6481), .Y(dp.rf._abc_6362_n6482) );
	NAND2X1 NAND2X1_4471 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6482), .Y(dp.rf._abc_6362_n6483) );
	NAND2X1 NAND2X1_4472 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6471), .B(dp.rf._abc_6362_n6483), .Y(dp.rf._abc_6362_n6484) );
	NAND2X1 NAND2X1_4473 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6484), .Y(dp.rf._abc_6362_n6485) );
	NAND2X1 NAND2X1_4474 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6485), .Y(dp.rf._abc_6362_n6486) );
	NAND2X1 NAND2X1_4475 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<11>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6487) );
	INVX1 INVX1_131 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<11>), .Y(dp.rf._abc_6362_n6488) );
	NOR2X1 NOR2X1_478 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6488), .Y(dp.rf._abc_6362_n6489) );
	NOR2X1 NOR2X1_479 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6489), .Y(dp.rf._abc_6362_n6490) );
	NAND2X1 NAND2X1_4476 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6487), .B(dp.rf._abc_6362_n6490), .Y(dp.rf._abc_6362_n6491) );
	NAND2X1 NAND2X1_4477 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<11>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6492) );
	INVX1 INVX1_132 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<11>), .Y(dp.rf._abc_6362_n6493) );
	NOR2X1 NOR2X1_480 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6493), .Y(dp.rf._abc_6362_n6494) );
	NOR2X1 NOR2X1_481 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6494), .Y(dp.rf._abc_6362_n6495) );
	NAND2X1 NAND2X1_4478 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6492), .B(dp.rf._abc_6362_n6495), .Y(dp.rf._abc_6362_n6496) );
	NAND2X1 NAND2X1_4479 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6491), .B(dp.rf._abc_6362_n6496), .Y(dp.rf._abc_6362_n6497) );
	NOR2X1 NOR2X1_482 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6497), .Y(dp.rf._abc_6362_n6498) );
	NAND2X1 NAND2X1_4480 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<11>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6499) );
	INVX1 INVX1_133 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<11>), .Y(dp.rf._abc_6362_n6500) );
	NOR2X1 NOR2X1_483 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6500), .Y(dp.rf._abc_6362_n6501) );
	NOR2X1 NOR2X1_484 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6501), .Y(dp.rf._abc_6362_n6502) );
	NAND2X1 NAND2X1_4481 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6499), .B(dp.rf._abc_6362_n6502), .Y(dp.rf._abc_6362_n6503) );
	NAND2X1 NAND2X1_4482 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<11>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6504) );
	INVX1 INVX1_134 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<11>), .Y(dp.rf._abc_6362_n6505) );
	NOR2X1 NOR2X1_485 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6505), .Y(dp.rf._abc_6362_n6506) );
	NOR2X1 NOR2X1_486 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6506), .Y(dp.rf._abc_6362_n6507) );
	NAND2X1 NAND2X1_4483 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6504), .B(dp.rf._abc_6362_n6507), .Y(dp.rf._abc_6362_n6508) );
	NAND2X1 NAND2X1_4484 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6503), .B(dp.rf._abc_6362_n6508), .Y(dp.rf._abc_6362_n6509) );
	NOR2X1 NOR2X1_487 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6509), .Y(dp.rf._abc_6362_n6510) );
	NOR2X1 NOR2X1_488 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6498), .B(dp.rf._abc_6362_n6510), .Y(dp.rf._abc_6362_n6511) );
	NOR2X1 NOR2X1_489 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6511), .Y(dp.rf._abc_6362_n6512) );
	NOR2X1 NOR2X1_490 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6486), .B(dp.rf._abc_6362_n6512), .Y(dp.rf._abc_6362_n6513) );
	NAND2X1 NAND2X1_4485 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<11>), .Y(dp.rf._abc_6362_n6514) );
	NAND2X1 NAND2X1_4486 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6514), .Y(dp.rf._abc_6362_n6515) );
	INVX1 INVX1_135 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<11>), .Y(dp.rf._abc_6362_n6516) );
	NOR2X1 NOR2X1_491 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6516), .Y(dp.rf._abc_6362_n6517) );
	NOR2X1 NOR2X1_492 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6515), .B(dp.rf._abc_6362_n6517), .Y(dp.rf._abc_6362_n6518) );
	NAND2X1 NAND2X1_4487 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<11>), .Y(dp.rf._abc_6362_n6519) );
	NAND2X1 NAND2X1_4488 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6519), .Y(dp.rf._abc_6362_n6520) );
	INVX1 INVX1_136 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<11>), .Y(dp.rf._abc_6362_n6521) );
	NOR2X1 NOR2X1_493 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6521), .Y(dp.rf._abc_6362_n6522) );
	NOR2X1 NOR2X1_494 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6520), .B(dp.rf._abc_6362_n6522), .Y(dp.rf._abc_6362_n6523) );
	OR2X2 OR2X2_47 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6518), .B(dp.rf._abc_6362_n6523), .Y(dp.rf._abc_6362_n6524) );
	NAND2X1 NAND2X1_4489 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6524), .Y(dp.rf._abc_6362_n6525) );
	NAND2X1 NAND2X1_4490 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<11>), .Y(dp.rf._abc_6362_n6526) );
	NAND2X1 NAND2X1_4491 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6526), .Y(dp.rf._abc_6362_n6527) );
	INVX1 INVX1_137 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<11>), .Y(dp.rf._abc_6362_n6528) );
	NOR2X1 NOR2X1_495 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6528), .Y(dp.rf._abc_6362_n6529) );
	NOR2X1 NOR2X1_496 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6527), .B(dp.rf._abc_6362_n6529), .Y(dp.rf._abc_6362_n6530) );
	NAND2X1 NAND2X1_4492 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<11>), .Y(dp.rf._abc_6362_n6531) );
	NAND2X1 NAND2X1_4493 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6531), .Y(dp.rf._abc_6362_n6532) );
	INVX1 INVX1_138 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<11>), .Y(dp.rf._abc_6362_n6533) );
	NOR2X1 NOR2X1_497 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6533), .Y(dp.rf._abc_6362_n6534) );
	NOR2X1 NOR2X1_498 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6532), .B(dp.rf._abc_6362_n6534), .Y(dp.rf._abc_6362_n6535) );
	OR2X2 OR2X2_48 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6530), .B(dp.rf._abc_6362_n6535), .Y(dp.rf._abc_6362_n6536) );
	NAND2X1 NAND2X1_4494 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6536), .Y(dp.rf._abc_6362_n6537) );
	AND2X2 AND2X2_169 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6537), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n6538) );
	NAND2X1 NAND2X1_4495 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6525), .B(dp.rf._abc_6362_n6538), .Y(dp.rf._abc_6362_n6539) );
	NAND2X1 NAND2X1_4496 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<11>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6540) );
	NAND2X1 NAND2X1_4497 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<11>), .Y(dp.rf._abc_6362_n6541) );
	AND2X2 AND2X2_170 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6541), .B(instr[22]), .Y(dp.rf._abc_6362_n6542) );
	NAND2X1 NAND2X1_4498 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6540), .B(dp.rf._abc_6362_n6542), .Y(dp.rf._abc_6362_n6543) );
	NAND2X1 NAND2X1_4499 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<11>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6544) );
	NAND2X1 NAND2X1_4500 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<11>), .Y(dp.rf._abc_6362_n6545) );
	AND2X2 AND2X2_171 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6545), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6546) );
	NAND2X1 NAND2X1_4501 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6544), .B(dp.rf._abc_6362_n6546), .Y(dp.rf._abc_6362_n6547) );
	NAND2X1 NAND2X1_4502 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6543), .B(dp.rf._abc_6362_n6547), .Y(dp.rf._abc_6362_n6548) );
	AND2X2 AND2X2_172 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6548), .B(instr[23]), .Y(dp.rf._abc_6362_n6549) );
	NAND2X1 NAND2X1_4503 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<11>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6550) );
	NAND2X1 NAND2X1_4504 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<11>), .Y(dp.rf._abc_6362_n6551) );
	AND2X2 AND2X2_173 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6551), .B(instr[22]), .Y(dp.rf._abc_6362_n6552) );
	NAND2X1 NAND2X1_4505 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6550), .B(dp.rf._abc_6362_n6552), .Y(dp.rf._abc_6362_n6553) );
	NAND2X1 NAND2X1_4506 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<11>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6554) );
	NAND2X1 NAND2X1_4507 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<11>), .Y(dp.rf._abc_6362_n6555) );
	AND2X2 AND2X2_174 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6555), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6556) );
	NAND2X1 NAND2X1_4508 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6554), .B(dp.rf._abc_6362_n6556), .Y(dp.rf._abc_6362_n6557) );
	NAND2X1 NAND2X1_4509 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6553), .B(dp.rf._abc_6362_n6557), .Y(dp.rf._abc_6362_n6558) );
	NAND2X1 NAND2X1_4510 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6558), .Y(dp.rf._abc_6362_n6559) );
	NAND2X1 NAND2X1_4511 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6559), .Y(dp.rf._abc_6362_n6560) );
	NOR2X1 NOR2X1_499 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6549), .B(dp.rf._abc_6362_n6560), .Y(dp.rf._abc_6362_n6561) );
	NOR2X1 NOR2X1_500 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6561), .Y(dp.rf._abc_6362_n6562) );
	NAND2X1 NAND2X1_4512 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6539), .B(dp.rf._abc_6362_n6562), .Y(dp.rf._abc_6362_n6563) );
	NAND2X1 NAND2X1_4513 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n6563), .Y(dp.rf._abc_6362_n6564) );
	NOR2X1 NOR2X1_501 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6513), .B(dp.rf._abc_6362_n6564), .Y(dp.srca_11_) );
	NAND2X1 NAND2X1_4514 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6566) );
	INVX1 INVX1_139 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<12>), .Y(dp.rf._abc_6362_n6567) );
	NOR2X1 NOR2X1_502 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6567), .Y(dp.rf._abc_6362_n6568) );
	NOR2X1 NOR2X1_503 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6568), .Y(dp.rf._abc_6362_n6569) );
	NAND2X1 NAND2X1_4515 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6566), .B(dp.rf._abc_6362_n6569), .Y(dp.rf._abc_6362_n6570) );
	NAND2X1 NAND2X1_4516 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6571) );
	INVX1 INVX1_140 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<12>), .Y(dp.rf._abc_6362_n6572) );
	NOR2X1 NOR2X1_504 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6572), .Y(dp.rf._abc_6362_n6573) );
	NOR2X1 NOR2X1_505 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6573), .Y(dp.rf._abc_6362_n6574) );
	NAND2X1 NAND2X1_4517 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6571), .B(dp.rf._abc_6362_n6574), .Y(dp.rf._abc_6362_n6575) );
	NAND2X1 NAND2X1_4518 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6570), .B(dp.rf._abc_6362_n6575), .Y(dp.rf._abc_6362_n6576) );
	NOR2X1 NOR2X1_506 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6576), .Y(dp.rf._abc_6362_n6577) );
	NAND2X1 NAND2X1_4519 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6578) );
	INVX1 INVX1_141 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<12>), .Y(dp.rf._abc_6362_n6579) );
	NOR2X1 NOR2X1_507 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6579), .Y(dp.rf._abc_6362_n6580) );
	NOR2X1 NOR2X1_508 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6580), .Y(dp.rf._abc_6362_n6581) );
	NAND2X1 NAND2X1_4520 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6578), .B(dp.rf._abc_6362_n6581), .Y(dp.rf._abc_6362_n6582) );
	NAND2X1 NAND2X1_4521 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6583) );
	INVX1 INVX1_142 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<12>), .Y(dp.rf._abc_6362_n6584) );
	NOR2X1 NOR2X1_509 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6584), .Y(dp.rf._abc_6362_n6585) );
	NOR2X1 NOR2X1_510 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6585), .Y(dp.rf._abc_6362_n6586) );
	NAND2X1 NAND2X1_4522 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6583), .B(dp.rf._abc_6362_n6586), .Y(dp.rf._abc_6362_n6587) );
	NAND2X1 NAND2X1_4523 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6582), .B(dp.rf._abc_6362_n6587), .Y(dp.rf._abc_6362_n6588) );
	NOR2X1 NOR2X1_511 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6588), .Y(dp.rf._abc_6362_n6589) );
	NOR2X1 NOR2X1_512 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6577), .B(dp.rf._abc_6362_n6589), .Y(dp.rf._abc_6362_n6590) );
	NOR2X1 NOR2X1_513 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6590), .Y(dp.rf._abc_6362_n6591) );
	NAND2X1 NAND2X1_4524 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<12>), .Y(dp.rf._abc_6362_n6592) );
	NAND2X1 NAND2X1_4525 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6592), .Y(dp.rf._abc_6362_n6593) );
	INVX1 INVX1_143 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<12>), .Y(dp.rf._abc_6362_n6594) );
	NOR2X1 NOR2X1_514 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6594), .Y(dp.rf._abc_6362_n6595) );
	NOR2X1 NOR2X1_515 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6593), .B(dp.rf._abc_6362_n6595), .Y(dp.rf._abc_6362_n6596) );
	NAND2X1 NAND2X1_4526 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<12>), .Y(dp.rf._abc_6362_n6597) );
	NAND2X1 NAND2X1_4527 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6597), .Y(dp.rf._abc_6362_n6598) );
	INVX1 INVX1_144 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<12>), .Y(dp.rf._abc_6362_n6599) );
	NOR2X1 NOR2X1_516 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6599), .Y(dp.rf._abc_6362_n6600) );
	NOR2X1 NOR2X1_517 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6598), .B(dp.rf._abc_6362_n6600), .Y(dp.rf._abc_6362_n6601) );
	OR2X2 OR2X2_49 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6596), .B(dp.rf._abc_6362_n6601), .Y(dp.rf._abc_6362_n6602) );
	NAND2X1 NAND2X1_4528 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6602), .Y(dp.rf._abc_6362_n6603) );
	NAND2X1 NAND2X1_4529 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<12>), .Y(dp.rf._abc_6362_n6604) );
	NAND2X1 NAND2X1_4530 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6604), .Y(dp.rf._abc_6362_n6605) );
	INVX1 INVX1_145 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<12>), .Y(dp.rf._abc_6362_n6606) );
	NOR2X1 NOR2X1_518 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6606), .Y(dp.rf._abc_6362_n6607) );
	NOR2X1 NOR2X1_519 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6605), .B(dp.rf._abc_6362_n6607), .Y(dp.rf._abc_6362_n6608) );
	NAND2X1 NAND2X1_4531 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<12>), .Y(dp.rf._abc_6362_n6609) );
	NAND2X1 NAND2X1_4532 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6609), .Y(dp.rf._abc_6362_n6610) );
	INVX1 INVX1_146 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<12>), .Y(dp.rf._abc_6362_n6611) );
	NOR2X1 NOR2X1_520 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6611), .Y(dp.rf._abc_6362_n6612) );
	NOR2X1 NOR2X1_521 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6610), .B(dp.rf._abc_6362_n6612), .Y(dp.rf._abc_6362_n6613) );
	OR2X2 OR2X2_50 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6608), .B(dp.rf._abc_6362_n6613), .Y(dp.rf._abc_6362_n6614) );
	NAND2X1 NAND2X1_4533 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6614), .Y(dp.rf._abc_6362_n6615) );
	AND2X2 AND2X2_175 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6615), .B(instr[24]), .Y(dp.rf._abc_6362_n6616) );
	NAND2X1 NAND2X1_4534 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6603), .B(dp.rf._abc_6362_n6616), .Y(dp.rf._abc_6362_n6617) );
	NAND2X1 NAND2X1_4535 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6617), .Y(dp.rf._abc_6362_n6618) );
	NOR2X1 NOR2X1_522 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6591), .B(dp.rf._abc_6362_n6618), .Y(dp.rf._abc_6362_n6619) );
	NAND2X1 NAND2X1_4536 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<12>), .Y(dp.rf._abc_6362_n6620) );
	NAND2X1 NAND2X1_4537 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6621) );
	NAND2X1 NAND2X1_4538 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6620), .B(dp.rf._abc_6362_n6621), .Y(dp.rf._abc_6362_n6622) );
	NAND2X1 NAND2X1_4539 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6622), .Y(dp.rf._abc_6362_n6623) );
	NAND2X1 NAND2X1_4540 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<12>), .Y(dp.rf._abc_6362_n6624) );
	NAND2X1 NAND2X1_4541 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6625) );
	NAND2X1 NAND2X1_4542 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6624), .B(dp.rf._abc_6362_n6625), .Y(dp.rf._abc_6362_n6626) );
	NAND2X1 NAND2X1_4543 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6626), .Y(dp.rf._abc_6362_n6627) );
	AND2X2 AND2X2_176 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6623), .B(dp.rf._abc_6362_n6627), .Y(dp.rf._abc_6362_n6628) );
	NAND2X1 NAND2X1_4544 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6628), .Y(dp.rf._abc_6362_n6629) );
	NAND2X1 NAND2X1_4545 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<12>), .Y(dp.rf._abc_6362_n6630) );
	NAND2X1 NAND2X1_4546 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6631) );
	NAND2X1 NAND2X1_4547 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6630), .B(dp.rf._abc_6362_n6631), .Y(dp.rf._abc_6362_n6632) );
	NAND2X1 NAND2X1_4548 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6632), .Y(dp.rf._abc_6362_n6633) );
	NAND2X1 NAND2X1_4549 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<12>), .Y(dp.rf._abc_6362_n6634) );
	NAND2X1 NAND2X1_4550 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6635) );
	NAND2X1 NAND2X1_4551 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6634), .B(dp.rf._abc_6362_n6635), .Y(dp.rf._abc_6362_n6636) );
	NAND2X1 NAND2X1_4552 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6636), .Y(dp.rf._abc_6362_n6637) );
	AND2X2 AND2X2_177 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6633), .B(dp.rf._abc_6362_n6637), .Y(dp.rf._abc_6362_n6638) );
	NAND2X1 NAND2X1_4553 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6638), .Y(dp.rf._abc_6362_n6639) );
	AND2X2 AND2X2_178 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6639), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n6640) );
	NAND2X1 NAND2X1_4554 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6629), .B(dp.rf._abc_6362_n6640), .Y(dp.rf._abc_6362_n6641) );
	NAND2X1 NAND2X1_4555 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6642) );
	NAND2X1 NAND2X1_4556 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<12>), .Y(dp.rf._abc_6362_n6643) );
	AND2X2 AND2X2_179 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6643), .B(instr[22]), .Y(dp.rf._abc_6362_n6644) );
	NAND2X1 NAND2X1_4557 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6642), .B(dp.rf._abc_6362_n6644), .Y(dp.rf._abc_6362_n6645) );
	NAND2X1 NAND2X1_4558 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6646) );
	NAND2X1 NAND2X1_4559 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<12>), .Y(dp.rf._abc_6362_n6647) );
	AND2X2 AND2X2_180 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6647), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6648) );
	NAND2X1 NAND2X1_4560 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6646), .B(dp.rf._abc_6362_n6648), .Y(dp.rf._abc_6362_n6649) );
	NAND2X1 NAND2X1_4561 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6645), .B(dp.rf._abc_6362_n6649), .Y(dp.rf._abc_6362_n6650) );
	AND2X2 AND2X2_181 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6650), .B(instr[23]), .Y(dp.rf._abc_6362_n6651) );
	NAND2X1 NAND2X1_4562 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6652) );
	NAND2X1 NAND2X1_4563 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<12>), .Y(dp.rf._abc_6362_n6653) );
	AND2X2 AND2X2_182 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6653), .B(instr[22]), .Y(dp.rf._abc_6362_n6654) );
	NAND2X1 NAND2X1_4564 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6652), .B(dp.rf._abc_6362_n6654), .Y(dp.rf._abc_6362_n6655) );
	NAND2X1 NAND2X1_4565 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<12>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6656) );
	NAND2X1 NAND2X1_4566 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<12>), .Y(dp.rf._abc_6362_n6657) );
	AND2X2 AND2X2_183 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6657), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6658) );
	NAND2X1 NAND2X1_4567 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6656), .B(dp.rf._abc_6362_n6658), .Y(dp.rf._abc_6362_n6659) );
	NAND2X1 NAND2X1_4568 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6655), .B(dp.rf._abc_6362_n6659), .Y(dp.rf._abc_6362_n6660) );
	NAND2X1 NAND2X1_4569 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6660), .Y(dp.rf._abc_6362_n6661) );
	NAND2X1 NAND2X1_4570 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6661), .Y(dp.rf._abc_6362_n6662) );
	NOR2X1 NOR2X1_523 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6651), .B(dp.rf._abc_6362_n6662), .Y(dp.rf._abc_6362_n6663) );
	NOR2X1 NOR2X1_524 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6663), .Y(dp.rf._abc_6362_n6664) );
	NAND2X1 NAND2X1_4571 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6641), .B(dp.rf._abc_6362_n6664), .Y(dp.rf._abc_6362_n6665) );
	NAND2X1 NAND2X1_4572 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n6665), .Y(dp.rf._abc_6362_n6666) );
	NOR2X1 NOR2X1_525 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6619), .B(dp.rf._abc_6362_n6666), .Y(dp.srca_12_) );
	NAND2X1 NAND2X1_4573 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<13>), .Y(dp.rf._abc_6362_n6668) );
	NAND2X1 NAND2X1_4574 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6668), .Y(dp.rf._abc_6362_n6669) );
	INVX1 INVX1_147 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<13>), .Y(dp.rf._abc_6362_n6670) );
	NOR2X1 NOR2X1_526 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6670), .Y(dp.rf._abc_6362_n6671) );
	NOR2X1 NOR2X1_527 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6669), .B(dp.rf._abc_6362_n6671), .Y(dp.rf._abc_6362_n6672) );
	NAND2X1 NAND2X1_4575 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<13>), .Y(dp.rf._abc_6362_n6673) );
	NAND2X1 NAND2X1_4576 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6673), .Y(dp.rf._abc_6362_n6674) );
	INVX1 INVX1_148 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<13>), .Y(dp.rf._abc_6362_n6675) );
	NOR2X1 NOR2X1_528 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6675), .Y(dp.rf._abc_6362_n6676) );
	NOR2X1 NOR2X1_529 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6674), .B(dp.rf._abc_6362_n6676), .Y(dp.rf._abc_6362_n6677) );
	NOR2X1 NOR2X1_530 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6672), .B(dp.rf._abc_6362_n6677), .Y(dp.rf._abc_6362_n6678) );
	NAND2X1 NAND2X1_4577 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6678), .Y(dp.rf._abc_6362_n6679) );
	NAND2X1 NAND2X1_4578 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<13>), .Y(dp.rf._abc_6362_n6680) );
	NAND2X1 NAND2X1_4579 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6680), .Y(dp.rf._abc_6362_n6681) );
	INVX1 INVX1_149 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<13>), .Y(dp.rf._abc_6362_n6682) );
	NOR2X1 NOR2X1_531 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6682), .Y(dp.rf._abc_6362_n6683) );
	NOR2X1 NOR2X1_532 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6681), .B(dp.rf._abc_6362_n6683), .Y(dp.rf._abc_6362_n6684) );
	NAND2X1 NAND2X1_4580 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<13>), .Y(dp.rf._abc_6362_n6685) );
	NAND2X1 NAND2X1_4581 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6685), .Y(dp.rf._abc_6362_n6686) );
	INVX1 INVX1_150 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<13>), .Y(dp.rf._abc_6362_n6687) );
	NOR2X1 NOR2X1_533 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6687), .Y(dp.rf._abc_6362_n6688) );
	NOR2X1 NOR2X1_534 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6686), .B(dp.rf._abc_6362_n6688), .Y(dp.rf._abc_6362_n6689) );
	NOR2X1 NOR2X1_535 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6684), .B(dp.rf._abc_6362_n6689), .Y(dp.rf._abc_6362_n6690) );
	NAND2X1 NAND2X1_4582 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6690), .Y(dp.rf._abc_6362_n6691) );
	NAND2X1 NAND2X1_4583 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6679), .B(dp.rf._abc_6362_n6691), .Y(dp.rf._abc_6362_n6692) );
	NAND2X1 NAND2X1_4584 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6692), .Y(dp.rf._abc_6362_n6693) );
	NAND2X1 NAND2X1_4585 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6693), .Y(dp.rf._abc_6362_n6694) );
	NAND2X1 NAND2X1_4586 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6695) );
	INVX1 INVX1_151 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<13>), .Y(dp.rf._abc_6362_n6696) );
	NOR2X1 NOR2X1_536 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6696), .Y(dp.rf._abc_6362_n6697) );
	NOR2X1 NOR2X1_537 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6697), .Y(dp.rf._abc_6362_n6698) );
	NAND2X1 NAND2X1_4587 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6695), .B(dp.rf._abc_6362_n6698), .Y(dp.rf._abc_6362_n6699) );
	NAND2X1 NAND2X1_4588 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6700) );
	INVX1 INVX1_152 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<13>), .Y(dp.rf._abc_6362_n6701) );
	NOR2X1 NOR2X1_538 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6701), .Y(dp.rf._abc_6362_n6702) );
	NOR2X1 NOR2X1_539 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6702), .Y(dp.rf._abc_6362_n6703) );
	NAND2X1 NAND2X1_4589 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6700), .B(dp.rf._abc_6362_n6703), .Y(dp.rf._abc_6362_n6704) );
	NAND2X1 NAND2X1_4590 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6699), .B(dp.rf._abc_6362_n6704), .Y(dp.rf._abc_6362_n6705) );
	NOR2X1 NOR2X1_540 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6705), .Y(dp.rf._abc_6362_n6706) );
	NAND2X1 NAND2X1_4591 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6707) );
	INVX1 INVX1_153 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<13>), .Y(dp.rf._abc_6362_n6708) );
	NOR2X1 NOR2X1_541 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6708), .Y(dp.rf._abc_6362_n6709) );
	NOR2X1 NOR2X1_542 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6709), .Y(dp.rf._abc_6362_n6710) );
	NAND2X1 NAND2X1_4592 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6707), .B(dp.rf._abc_6362_n6710), .Y(dp.rf._abc_6362_n6711) );
	NAND2X1 NAND2X1_4593 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6712) );
	INVX1 INVX1_154 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<13>), .Y(dp.rf._abc_6362_n6713) );
	NOR2X1 NOR2X1_543 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6713), .Y(dp.rf._abc_6362_n6714) );
	NOR2X1 NOR2X1_544 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6714), .Y(dp.rf._abc_6362_n6715) );
	NAND2X1 NAND2X1_4594 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6712), .B(dp.rf._abc_6362_n6715), .Y(dp.rf._abc_6362_n6716) );
	NAND2X1 NAND2X1_4595 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6711), .B(dp.rf._abc_6362_n6716), .Y(dp.rf._abc_6362_n6717) );
	NOR2X1 NOR2X1_545 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6717), .Y(dp.rf._abc_6362_n6718) );
	NOR2X1 NOR2X1_546 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6706), .B(dp.rf._abc_6362_n6718), .Y(dp.rf._abc_6362_n6719) );
	NOR2X1 NOR2X1_547 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6719), .Y(dp.rf._abc_6362_n6720) );
	NOR2X1 NOR2X1_548 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6694), .B(dp.rf._abc_6362_n6720), .Y(dp.rf._abc_6362_n6721) );
	NAND2X1 NAND2X1_4596 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<13>), .Y(dp.rf._abc_6362_n6722) );
	NAND2X1 NAND2X1_4597 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6723) );
	NAND2X1 NAND2X1_4598 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6722), .B(dp.rf._abc_6362_n6723), .Y(dp.rf._abc_6362_n6724) );
	NAND2X1 NAND2X1_4599 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6724), .Y(dp.rf._abc_6362_n6725) );
	NAND2X1 NAND2X1_4600 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<13>), .Y(dp.rf._abc_6362_n6726) );
	NAND2X1 NAND2X1_4601 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6727) );
	NAND2X1 NAND2X1_4602 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6726), .B(dp.rf._abc_6362_n6727), .Y(dp.rf._abc_6362_n6728) );
	NAND2X1 NAND2X1_4603 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6728), .Y(dp.rf._abc_6362_n6729) );
	AND2X2 AND2X2_184 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6725), .B(dp.rf._abc_6362_n6729), .Y(dp.rf._abc_6362_n6730) );
	NAND2X1 NAND2X1_4604 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6730), .Y(dp.rf._abc_6362_n6731) );
	NAND2X1 NAND2X1_4605 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<13>), .Y(dp.rf._abc_6362_n6732) );
	NAND2X1 NAND2X1_4606 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6733) );
	NAND2X1 NAND2X1_4607 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6732), .B(dp.rf._abc_6362_n6733), .Y(dp.rf._abc_6362_n6734) );
	NAND2X1 NAND2X1_4608 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6734), .Y(dp.rf._abc_6362_n6735) );
	NAND2X1 NAND2X1_4609 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<13>), .Y(dp.rf._abc_6362_n6736) );
	NAND2X1 NAND2X1_4610 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6737) );
	NAND2X1 NAND2X1_4611 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6736), .B(dp.rf._abc_6362_n6737), .Y(dp.rf._abc_6362_n6738) );
	NAND2X1 NAND2X1_4612 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6738), .Y(dp.rf._abc_6362_n6739) );
	AND2X2 AND2X2_185 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6735), .B(dp.rf._abc_6362_n6739), .Y(dp.rf._abc_6362_n6740) );
	NAND2X1 NAND2X1_4613 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6740), .Y(dp.rf._abc_6362_n6741) );
	AND2X2 AND2X2_186 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6741), .B(instr[24]), .Y(dp.rf._abc_6362_n6742) );
	NAND2X1 NAND2X1_4614 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6731), .B(dp.rf._abc_6362_n6742), .Y(dp.rf._abc_6362_n6743) );
	NAND2X1 NAND2X1_4615 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6744) );
	NAND2X1 NAND2X1_4616 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<13>), .Y(dp.rf._abc_6362_n6745) );
	AND2X2 AND2X2_187 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6745), .B(instr[22]), .Y(dp.rf._abc_6362_n6746) );
	NAND2X1 NAND2X1_4617 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6744), .B(dp.rf._abc_6362_n6746), .Y(dp.rf._abc_6362_n6747) );
	NAND2X1 NAND2X1_4618 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6748) );
	NAND2X1 NAND2X1_4619 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<13>), .Y(dp.rf._abc_6362_n6749) );
	AND2X2 AND2X2_188 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6749), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6750) );
	NAND2X1 NAND2X1_4620 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6748), .B(dp.rf._abc_6362_n6750), .Y(dp.rf._abc_6362_n6751) );
	NAND2X1 NAND2X1_4621 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6747), .B(dp.rf._abc_6362_n6751), .Y(dp.rf._abc_6362_n6752) );
	AND2X2 AND2X2_189 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6752), .B(instr[23]), .Y(dp.rf._abc_6362_n6753) );
	NAND2X1 NAND2X1_4622 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6754) );
	NAND2X1 NAND2X1_4623 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<13>), .Y(dp.rf._abc_6362_n6755) );
	AND2X2 AND2X2_190 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6755), .B(instr[22]), .Y(dp.rf._abc_6362_n6756) );
	NAND2X1 NAND2X1_4624 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6754), .B(dp.rf._abc_6362_n6756), .Y(dp.rf._abc_6362_n6757) );
	NAND2X1 NAND2X1_4625 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<13>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6758) );
	NAND2X1 NAND2X1_4626 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<13>), .Y(dp.rf._abc_6362_n6759) );
	AND2X2 AND2X2_191 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6759), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6760) );
	NAND2X1 NAND2X1_4627 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6758), .B(dp.rf._abc_6362_n6760), .Y(dp.rf._abc_6362_n6761) );
	NAND2X1 NAND2X1_4628 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6757), .B(dp.rf._abc_6362_n6761), .Y(dp.rf._abc_6362_n6762) );
	NAND2X1 NAND2X1_4629 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6762), .Y(dp.rf._abc_6362_n6763) );
	NAND2X1 NAND2X1_4630 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n6763), .Y(dp.rf._abc_6362_n6764) );
	NOR2X1 NOR2X1_549 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6753), .B(dp.rf._abc_6362_n6764), .Y(dp.rf._abc_6362_n6765) );
	NOR2X1 NOR2X1_550 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6765), .Y(dp.rf._abc_6362_n6766) );
	NAND2X1 NAND2X1_4631 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6743), .B(dp.rf._abc_6362_n6766), .Y(dp.rf._abc_6362_n6767) );
	NAND2X1 NAND2X1_4632 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n6767), .Y(dp.rf._abc_6362_n6768) );
	NOR2X1 NOR2X1_551 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6721), .B(dp.rf._abc_6362_n6768), .Y(dp.srca_13_) );
	NAND2X1 NAND2X1_4633 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<14>), .Y(dp.rf._abc_6362_n6770) );
	NAND2X1 NAND2X1_4634 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6770), .Y(dp.rf._abc_6362_n6771) );
	INVX1 INVX1_155 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<14>), .Y(dp.rf._abc_6362_n6772) );
	NOR2X1 NOR2X1_552 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6772), .Y(dp.rf._abc_6362_n6773) );
	NOR2X1 NOR2X1_553 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6771), .B(dp.rf._abc_6362_n6773), .Y(dp.rf._abc_6362_n6774) );
	NAND2X1 NAND2X1_4635 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<14>), .Y(dp.rf._abc_6362_n6775) );
	NAND2X1 NAND2X1_4636 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6775), .Y(dp.rf._abc_6362_n6776) );
	INVX1 INVX1_156 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<14>), .Y(dp.rf._abc_6362_n6777) );
	NOR2X1 NOR2X1_554 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6777), .Y(dp.rf._abc_6362_n6778) );
	NOR2X1 NOR2X1_555 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6776), .B(dp.rf._abc_6362_n6778), .Y(dp.rf._abc_6362_n6779) );
	NOR2X1 NOR2X1_556 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6774), .B(dp.rf._abc_6362_n6779), .Y(dp.rf._abc_6362_n6780) );
	NAND2X1 NAND2X1_4637 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6780), .Y(dp.rf._abc_6362_n6781) );
	NAND2X1 NAND2X1_4638 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<14>), .Y(dp.rf._abc_6362_n6782) );
	NAND2X1 NAND2X1_4639 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6782), .Y(dp.rf._abc_6362_n6783) );
	INVX1 INVX1_157 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<14>), .Y(dp.rf._abc_6362_n6784) );
	NOR2X1 NOR2X1_557 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6784), .Y(dp.rf._abc_6362_n6785) );
	NOR2X1 NOR2X1_558 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6783), .B(dp.rf._abc_6362_n6785), .Y(dp.rf._abc_6362_n6786) );
	NAND2X1 NAND2X1_4640 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<14>), .Y(dp.rf._abc_6362_n6787) );
	NAND2X1 NAND2X1_4641 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6787), .Y(dp.rf._abc_6362_n6788) );
	INVX1 INVX1_158 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<14>), .Y(dp.rf._abc_6362_n6789) );
	NOR2X1 NOR2X1_559 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6789), .Y(dp.rf._abc_6362_n6790) );
	NOR2X1 NOR2X1_560 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6788), .B(dp.rf._abc_6362_n6790), .Y(dp.rf._abc_6362_n6791) );
	NOR2X1 NOR2X1_561 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6786), .B(dp.rf._abc_6362_n6791), .Y(dp.rf._abc_6362_n6792) );
	NAND2X1 NAND2X1_4642 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6792), .Y(dp.rf._abc_6362_n6793) );
	NAND2X1 NAND2X1_4643 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6781), .B(dp.rf._abc_6362_n6793), .Y(dp.rf._abc_6362_n6794) );
	NAND2X1 NAND2X1_4644 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6794), .Y(dp.rf._abc_6362_n6795) );
	NAND2X1 NAND2X1_4645 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6795), .Y(dp.rf._abc_6362_n6796) );
	NAND2X1 NAND2X1_4646 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6797) );
	INVX1 INVX1_159 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<14>), .Y(dp.rf._abc_6362_n6798) );
	NOR2X1 NOR2X1_562 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6798), .Y(dp.rf._abc_6362_n6799) );
	NOR2X1 NOR2X1_563 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6799), .Y(dp.rf._abc_6362_n6800) );
	NAND2X1 NAND2X1_4647 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6797), .B(dp.rf._abc_6362_n6800), .Y(dp.rf._abc_6362_n6801) );
	NAND2X1 NAND2X1_4648 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6802) );
	INVX1 INVX1_160 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<14>), .Y(dp.rf._abc_6362_n6803) );
	NOR2X1 NOR2X1_564 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6803), .Y(dp.rf._abc_6362_n6804) );
	NOR2X1 NOR2X1_565 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6804), .Y(dp.rf._abc_6362_n6805) );
	NAND2X1 NAND2X1_4649 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6802), .B(dp.rf._abc_6362_n6805), .Y(dp.rf._abc_6362_n6806) );
	NAND2X1 NAND2X1_4650 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6801), .B(dp.rf._abc_6362_n6806), .Y(dp.rf._abc_6362_n6807) );
	NOR2X1 NOR2X1_566 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6807), .Y(dp.rf._abc_6362_n6808) );
	NAND2X1 NAND2X1_4651 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6809) );
	INVX1 INVX1_161 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<14>), .Y(dp.rf._abc_6362_n6810) );
	NOR2X1 NOR2X1_567 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6810), .Y(dp.rf._abc_6362_n6811) );
	NOR2X1 NOR2X1_568 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6811), .Y(dp.rf._abc_6362_n6812) );
	NAND2X1 NAND2X1_4652 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6809), .B(dp.rf._abc_6362_n6812), .Y(dp.rf._abc_6362_n6813) );
	NAND2X1 NAND2X1_4653 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6814) );
	INVX1 INVX1_162 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<14>), .Y(dp.rf._abc_6362_n6815) );
	NOR2X1 NOR2X1_569 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n6815), .Y(dp.rf._abc_6362_n6816) );
	NOR2X1 NOR2X1_570 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6816), .Y(dp.rf._abc_6362_n6817) );
	NAND2X1 NAND2X1_4654 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6814), .B(dp.rf._abc_6362_n6817), .Y(dp.rf._abc_6362_n6818) );
	NAND2X1 NAND2X1_4655 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6813), .B(dp.rf._abc_6362_n6818), .Y(dp.rf._abc_6362_n6819) );
	NOR2X1 NOR2X1_571 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6819), .Y(dp.rf._abc_6362_n6820) );
	NOR2X1 NOR2X1_572 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6808), .B(dp.rf._abc_6362_n6820), .Y(dp.rf._abc_6362_n6821) );
	NOR2X1 NOR2X1_573 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6821), .Y(dp.rf._abc_6362_n6822) );
	NOR2X1 NOR2X1_574 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6796), .B(dp.rf._abc_6362_n6822), .Y(dp.rf._abc_6362_n6823) );
	NAND2X1 NAND2X1_4656 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<14>), .Y(dp.rf._abc_6362_n6824) );
	NAND2X1 NAND2X1_4657 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6825) );
	NAND2X1 NAND2X1_4658 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6824), .B(dp.rf._abc_6362_n6825), .Y(dp.rf._abc_6362_n6826) );
	NAND2X1 NAND2X1_4659 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6826), .Y(dp.rf._abc_6362_n6827) );
	NAND2X1 NAND2X1_4660 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<14>), .Y(dp.rf._abc_6362_n6828) );
	NAND2X1 NAND2X1_4661 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6829) );
	NAND2X1 NAND2X1_4662 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6828), .B(dp.rf._abc_6362_n6829), .Y(dp.rf._abc_6362_n6830) );
	NAND2X1 NAND2X1_4663 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6830), .Y(dp.rf._abc_6362_n6831) );
	AND2X2 AND2X2_192 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6827), .B(dp.rf._abc_6362_n6831), .Y(dp.rf._abc_6362_n6832) );
	NAND2X1 NAND2X1_4664 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6832), .Y(dp.rf._abc_6362_n6833) );
	NAND2X1 NAND2X1_4665 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<14>), .Y(dp.rf._abc_6362_n6834) );
	NAND2X1 NAND2X1_4666 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6835) );
	NAND2X1 NAND2X1_4667 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6834), .B(dp.rf._abc_6362_n6835), .Y(dp.rf._abc_6362_n6836) );
	NAND2X1 NAND2X1_4668 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6836), .Y(dp.rf._abc_6362_n6837) );
	NAND2X1 NAND2X1_4669 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<14>), .Y(dp.rf._abc_6362_n6838) );
	NAND2X1 NAND2X1_4670 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6839) );
	NAND2X1 NAND2X1_4671 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6838), .B(dp.rf._abc_6362_n6839), .Y(dp.rf._abc_6362_n6840) );
	NAND2X1 NAND2X1_4672 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6840), .Y(dp.rf._abc_6362_n6841) );
	AND2X2 AND2X2_193 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6837), .B(dp.rf._abc_6362_n6841), .Y(dp.rf._abc_6362_n6842) );
	NAND2X1 NAND2X1_4673 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6842), .Y(dp.rf._abc_6362_n6843) );
	AND2X2 AND2X2_194 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6843), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n6844) );
	NAND2X1 NAND2X1_4674 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6833), .B(dp.rf._abc_6362_n6844), .Y(dp.rf._abc_6362_n6845) );
	NAND2X1 NAND2X1_4675 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6846) );
	NAND2X1 NAND2X1_4676 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<14>), .Y(dp.rf._abc_6362_n6847) );
	AND2X2 AND2X2_195 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6847), .B(instr[22]), .Y(dp.rf._abc_6362_n6848) );
	NAND2X1 NAND2X1_4677 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6846), .B(dp.rf._abc_6362_n6848), .Y(dp.rf._abc_6362_n6849) );
	NAND2X1 NAND2X1_4678 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6850) );
	NAND2X1 NAND2X1_4679 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<14>), .Y(dp.rf._abc_6362_n6851) );
	AND2X2 AND2X2_196 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6851), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6852) );
	NAND2X1 NAND2X1_4680 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6850), .B(dp.rf._abc_6362_n6852), .Y(dp.rf._abc_6362_n6853) );
	NAND2X1 NAND2X1_4681 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6849), .B(dp.rf._abc_6362_n6853), .Y(dp.rf._abc_6362_n6854) );
	AND2X2 AND2X2_197 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6854), .B(instr[23]), .Y(dp.rf._abc_6362_n6855) );
	NAND2X1 NAND2X1_4682 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6856) );
	NAND2X1 NAND2X1_4683 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<14>), .Y(dp.rf._abc_6362_n6857) );
	AND2X2 AND2X2_198 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6857), .B(instr[22]), .Y(dp.rf._abc_6362_n6858) );
	NAND2X1 NAND2X1_4684 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6856), .B(dp.rf._abc_6362_n6858), .Y(dp.rf._abc_6362_n6859) );
	NAND2X1 NAND2X1_4685 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<14>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6860) );
	NAND2X1 NAND2X1_4686 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<14>), .Y(dp.rf._abc_6362_n6861) );
	AND2X2 AND2X2_199 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6861), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6862) );
	NAND2X1 NAND2X1_4687 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6860), .B(dp.rf._abc_6362_n6862), .Y(dp.rf._abc_6362_n6863) );
	NAND2X1 NAND2X1_4688 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6859), .B(dp.rf._abc_6362_n6863), .Y(dp.rf._abc_6362_n6864) );
	NAND2X1 NAND2X1_4689 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6864), .Y(dp.rf._abc_6362_n6865) );
	NAND2X1 NAND2X1_4690 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6865), .Y(dp.rf._abc_6362_n6866) );
	NOR2X1 NOR2X1_575 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6855), .B(dp.rf._abc_6362_n6866), .Y(dp.rf._abc_6362_n6867) );
	NOR2X1 NOR2X1_576 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6867), .Y(dp.rf._abc_6362_n6868) );
	NAND2X1 NAND2X1_4691 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6845), .B(dp.rf._abc_6362_n6868), .Y(dp.rf._abc_6362_n6869) );
	NAND2X1 NAND2X1_4692 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n6869), .Y(dp.rf._abc_6362_n6870) );
	NOR2X1 NOR2X1_577 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6823), .B(dp.rf._abc_6362_n6870), .Y(dp.srca_14_) );
	NAND2X1 NAND2X1_4693 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<15>), .Y(dp.rf._abc_6362_n6872) );
	NAND2X1 NAND2X1_4694 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6873) );
	NAND2X1 NAND2X1_4695 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6872), .B(dp.rf._abc_6362_n6873), .Y(dp.rf._abc_6362_n6874) );
	NAND2X1 NAND2X1_4696 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6874), .Y(dp.rf._abc_6362_n6875) );
	NAND2X1 NAND2X1_4697 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<15>), .Y(dp.rf._abc_6362_n6876) );
	NAND2X1 NAND2X1_4698 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6877) );
	NAND2X1 NAND2X1_4699 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6876), .B(dp.rf._abc_6362_n6877), .Y(dp.rf._abc_6362_n6878) );
	NAND2X1 NAND2X1_4700 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6878), .Y(dp.rf._abc_6362_n6879) );
	NAND2X1 NAND2X1_4701 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6875), .B(dp.rf._abc_6362_n6879), .Y(dp.rf._abc_6362_n6880) );
	NOR2X1 NOR2X1_578 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6880), .Y(dp.rf._abc_6362_n6881) );
	NAND2X1 NAND2X1_4702 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<15>), .Y(dp.rf._abc_6362_n6882) );
	NAND2X1 NAND2X1_4703 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6883) );
	NAND2X1 NAND2X1_4704 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6882), .B(dp.rf._abc_6362_n6883), .Y(dp.rf._abc_6362_n6884) );
	NAND2X1 NAND2X1_4705 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6884), .Y(dp.rf._abc_6362_n6885) );
	NAND2X1 NAND2X1_4706 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<15>), .Y(dp.rf._abc_6362_n6886) );
	NAND2X1 NAND2X1_4707 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6887) );
	NAND2X1 NAND2X1_4708 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6886), .B(dp.rf._abc_6362_n6887), .Y(dp.rf._abc_6362_n6888) );
	NAND2X1 NAND2X1_4709 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6888), .Y(dp.rf._abc_6362_n6889) );
	AND2X2 AND2X2_200 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6885), .B(dp.rf._abc_6362_n6889), .Y(dp.rf._abc_6362_n6890) );
	NAND2X1 NAND2X1_4710 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6890), .Y(dp.rf._abc_6362_n6891) );
	NAND2X1 NAND2X1_4711 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n6891), .Y(dp.rf._abc_6362_n6892) );
	NOR2X1 NOR2X1_579 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6881), .B(dp.rf._abc_6362_n6892), .Y(dp.rf._abc_6362_n6893) );
	NAND2X1 NAND2X1_4712 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<15>), .Y(dp.rf._abc_6362_n6894) );
	NAND2X1 NAND2X1_4713 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6895) );
	NAND2X1 NAND2X1_4714 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6894), .B(dp.rf._abc_6362_n6895), .Y(dp.rf._abc_6362_n6896) );
	NAND2X1 NAND2X1_4715 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6896), .Y(dp.rf._abc_6362_n6897) );
	NAND2X1 NAND2X1_4716 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<15>), .Y(dp.rf._abc_6362_n6898) );
	NAND2X1 NAND2X1_4717 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6899) );
	NAND2X1 NAND2X1_4718 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6898), .B(dp.rf._abc_6362_n6899), .Y(dp.rf._abc_6362_n6900) );
	NAND2X1 NAND2X1_4719 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6900), .Y(dp.rf._abc_6362_n6901) );
	AND2X2 AND2X2_201 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6897), .B(dp.rf._abc_6362_n6901), .Y(dp.rf._abc_6362_n6902) );
	NAND2X1 NAND2X1_4720 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6902), .Y(dp.rf._abc_6362_n6903) );
	NAND2X1 NAND2X1_4721 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<15>), .Y(dp.rf._abc_6362_n6904) );
	NAND2X1 NAND2X1_4722 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6904), .Y(dp.rf._abc_6362_n6905) );
	AND2X2 AND2X2_202 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf.rf_10_<15>), .Y(dp.rf._abc_6362_n6906) );
	NOR2X1 NOR2X1_580 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6905), .B(dp.rf._abc_6362_n6906), .Y(dp.rf._abc_6362_n6907) );
	NAND2X1 NAND2X1_4723 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<15>), .Y(dp.rf._abc_6362_n6908) );
	NAND2X1 NAND2X1_4724 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6908), .Y(dp.rf._abc_6362_n6909) );
	INVX1 INVX1_163 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<15>), .Y(dp.rf._abc_6362_n6910) );
	NOR2X1 NOR2X1_581 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n6910), .Y(dp.rf._abc_6362_n6911) );
	NOR2X1 NOR2X1_582 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6909), .B(dp.rf._abc_6362_n6911), .Y(dp.rf._abc_6362_n6912) );
	OR2X2 OR2X2_51 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6907), .B(dp.rf._abc_6362_n6912), .Y(dp.rf._abc_6362_n6913) );
	NAND2X1 NAND2X1_4725 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6913), .Y(dp.rf._abc_6362_n6914) );
	AND2X2 AND2X2_203 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6914), .B(instr[24]), .Y(dp.rf._abc_6362_n6915) );
	NAND2X1 NAND2X1_4726 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6903), .B(dp.rf._abc_6362_n6915), .Y(dp.rf._abc_6362_n6916) );
	NAND2X1 NAND2X1_4727 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6916), .Y(dp.rf._abc_6362_n6917) );
	NOR2X1 NOR2X1_583 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6893), .B(dp.rf._abc_6362_n6917), .Y(dp.rf._abc_6362_n6918) );
	NAND2X1 NAND2X1_4728 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<15>), .Y(dp.rf._abc_6362_n6919) );
	NAND2X1 NAND2X1_4729 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6920) );
	NAND2X1 NAND2X1_4730 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6919), .B(dp.rf._abc_6362_n6920), .Y(dp.rf._abc_6362_n6921) );
	NAND2X1 NAND2X1_4731 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6921), .Y(dp.rf._abc_6362_n6922) );
	NAND2X1 NAND2X1_4732 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<15>), .Y(dp.rf._abc_6362_n6923) );
	NAND2X1 NAND2X1_4733 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6924) );
	NAND2X1 NAND2X1_4734 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6923), .B(dp.rf._abc_6362_n6924), .Y(dp.rf._abc_6362_n6925) );
	NAND2X1 NAND2X1_4735 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6925), .Y(dp.rf._abc_6362_n6926) );
	AND2X2 AND2X2_204 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6922), .B(dp.rf._abc_6362_n6926), .Y(dp.rf._abc_6362_n6927) );
	NAND2X1 NAND2X1_4736 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6927), .Y(dp.rf._abc_6362_n6928) );
	NAND2X1 NAND2X1_4737 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<15>), .Y(dp.rf._abc_6362_n6929) );
	NAND2X1 NAND2X1_4738 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6930) );
	NAND2X1 NAND2X1_4739 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6929), .B(dp.rf._abc_6362_n6930), .Y(dp.rf._abc_6362_n6931) );
	NAND2X1 NAND2X1_4740 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6931), .Y(dp.rf._abc_6362_n6932) );
	NAND2X1 NAND2X1_4741 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<15>), .Y(dp.rf._abc_6362_n6933) );
	NAND2X1 NAND2X1_4742 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6934) );
	NAND2X1 NAND2X1_4743 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6933), .B(dp.rf._abc_6362_n6934), .Y(dp.rf._abc_6362_n6935) );
	NAND2X1 NAND2X1_4744 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6935), .Y(dp.rf._abc_6362_n6936) );
	AND2X2 AND2X2_205 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6932), .B(dp.rf._abc_6362_n6936), .Y(dp.rf._abc_6362_n6937) );
	NAND2X1 NAND2X1_4745 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6937), .Y(dp.rf._abc_6362_n6938) );
	AND2X2 AND2X2_206 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6938), .B(instr[24]), .Y(dp.rf._abc_6362_n6939) );
	NAND2X1 NAND2X1_4746 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6928), .B(dp.rf._abc_6362_n6939), .Y(dp.rf._abc_6362_n6940) );
	NAND2X1 NAND2X1_4747 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6941) );
	NAND2X1 NAND2X1_4748 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<15>), .Y(dp.rf._abc_6362_n6942) );
	AND2X2 AND2X2_207 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6942), .B(instr[22]), .Y(dp.rf._abc_6362_n6943) );
	NAND2X1 NAND2X1_4749 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6941), .B(dp.rf._abc_6362_n6943), .Y(dp.rf._abc_6362_n6944) );
	NAND2X1 NAND2X1_4750 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6945) );
	NAND2X1 NAND2X1_4751 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<15>), .Y(dp.rf._abc_6362_n6946) );
	AND2X2 AND2X2_208 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6946), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6947) );
	NAND2X1 NAND2X1_4752 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6945), .B(dp.rf._abc_6362_n6947), .Y(dp.rf._abc_6362_n6948) );
	NAND2X1 NAND2X1_4753 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6944), .B(dp.rf._abc_6362_n6948), .Y(dp.rf._abc_6362_n6949) );
	AND2X2 AND2X2_209 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6949), .B(instr[23]), .Y(dp.rf._abc_6362_n6950) );
	NAND2X1 NAND2X1_4754 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6951) );
	NAND2X1 NAND2X1_4755 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<15>), .Y(dp.rf._abc_6362_n6952) );
	AND2X2 AND2X2_210 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6952), .B(instr[22]), .Y(dp.rf._abc_6362_n6953) );
	NAND2X1 NAND2X1_4756 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6951), .B(dp.rf._abc_6362_n6953), .Y(dp.rf._abc_6362_n6954) );
	NAND2X1 NAND2X1_4757 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<15>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6955) );
	NAND2X1 NAND2X1_4758 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<15>), .Y(dp.rf._abc_6362_n6956) );
	AND2X2 AND2X2_211 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6956), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n6957) );
	NAND2X1 NAND2X1_4759 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6955), .B(dp.rf._abc_6362_n6957), .Y(dp.rf._abc_6362_n6958) );
	NAND2X1 NAND2X1_4760 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6954), .B(dp.rf._abc_6362_n6958), .Y(dp.rf._abc_6362_n6959) );
	NAND2X1 NAND2X1_4761 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n6959), .Y(dp.rf._abc_6362_n6960) );
	NAND2X1 NAND2X1_4762 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n6960), .Y(dp.rf._abc_6362_n6961) );
	NOR2X1 NOR2X1_584 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6950), .B(dp.rf._abc_6362_n6961), .Y(dp.rf._abc_6362_n6962) );
	NOR2X1 NOR2X1_585 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n6962), .Y(dp.rf._abc_6362_n6963) );
	NAND2X1 NAND2X1_4763 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6940), .B(dp.rf._abc_6362_n6963), .Y(dp.rf._abc_6362_n6964) );
	NAND2X1 NAND2X1_4764 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n6964), .Y(dp.rf._abc_6362_n6965) );
	NOR2X1 NOR2X1_586 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6918), .B(dp.rf._abc_6362_n6965), .Y(dp.srca_15_) );
	NAND2X1 NAND2X1_4765 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<16>), .Y(dp.rf._abc_6362_n6967) );
	NAND2X1 NAND2X1_4766 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<16>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6968) );
	NAND2X1 NAND2X1_4767 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6967), .B(dp.rf._abc_6362_n6968), .Y(dp.rf._abc_6362_n6969) );
	NAND2X1 NAND2X1_4768 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6969), .Y(dp.rf._abc_6362_n6970) );
	NAND2X1 NAND2X1_4769 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<16>), .Y(dp.rf._abc_6362_n6971) );
	NAND2X1 NAND2X1_4770 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<16>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6972) );
	NAND2X1 NAND2X1_4771 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6971), .B(dp.rf._abc_6362_n6972), .Y(dp.rf._abc_6362_n6973) );
	NAND2X1 NAND2X1_4772 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6973), .Y(dp.rf._abc_6362_n6974) );
	NAND2X1 NAND2X1_4773 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6970), .B(dp.rf._abc_6362_n6974), .Y(dp.rf._abc_6362_n6975) );
	NOR2X1 NOR2X1_587 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6975), .Y(dp.rf._abc_6362_n6976) );
	NAND2X1 NAND2X1_4774 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<16>), .Y(dp.rf._abc_6362_n6977) );
	NAND2X1 NAND2X1_4775 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<16>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6978) );
	NAND2X1 NAND2X1_4776 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6977), .B(dp.rf._abc_6362_n6978), .Y(dp.rf._abc_6362_n6979) );
	NAND2X1 NAND2X1_4777 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6979), .Y(dp.rf._abc_6362_n6980) );
	NAND2X1 NAND2X1_4778 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<16>), .Y(dp.rf._abc_6362_n6981) );
	NAND2X1 NAND2X1_4779 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<16>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6982) );
	NAND2X1 NAND2X1_4780 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6981), .B(dp.rf._abc_6362_n6982), .Y(dp.rf._abc_6362_n6983) );
	NAND2X1 NAND2X1_4781 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6983), .Y(dp.rf._abc_6362_n6984) );
	AND2X2 AND2X2_212 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6980), .B(dp.rf._abc_6362_n6984), .Y(dp.rf._abc_6362_n6985) );
	NAND2X1 NAND2X1_4782 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6985), .Y(dp.rf._abc_6362_n6986) );
	NAND2X1 NAND2X1_4783 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n6986), .Y(dp.rf._abc_6362_n6987) );
	NOR2X1 NOR2X1_588 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6976), .B(dp.rf._abc_6362_n6987), .Y(dp.rf._abc_6362_n6988) );
	NAND2X1 NAND2X1_4784 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<16>), .Y(dp.rf._abc_6362_n6989) );
	NAND2X1 NAND2X1_4785 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<16>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6990) );
	NAND2X1 NAND2X1_4786 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6989), .B(dp.rf._abc_6362_n6990), .Y(dp.rf._abc_6362_n6991) );
	NAND2X1 NAND2X1_4787 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n6991), .Y(dp.rf._abc_6362_n6992) );
	NAND2X1 NAND2X1_4788 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<16>), .Y(dp.rf._abc_6362_n6993) );
	NAND2X1 NAND2X1_4789 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<16>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n6994) );
	NAND2X1 NAND2X1_4790 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6993), .B(dp.rf._abc_6362_n6994), .Y(dp.rf._abc_6362_n6995) );
	NAND2X1 NAND2X1_4791 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6995), .Y(dp.rf._abc_6362_n6996) );
	AND2X2 AND2X2_213 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6992), .B(dp.rf._abc_6362_n6996), .Y(dp.rf._abc_6362_n6997) );
	NAND2X1 NAND2X1_4792 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n6997), .Y(dp.rf._abc_6362_n6998) );
	NAND2X1 NAND2X1_4793 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<16>), .Y(dp.rf._abc_6362_n6999) );
	NAND2X1 NAND2X1_4794 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n6999), .Y(dp.rf._abc_6362_n7000) );
	AND2X2 AND2X2_214 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf.rf_2_<16>), .Y(dp.rf._abc_6362_n7001) );
	NOR2X1 NOR2X1_589 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7000), .B(dp.rf._abc_6362_n7001), .Y(dp.rf._abc_6362_n7002) );
	NAND2X1 NAND2X1_4795 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<16>), .Y(dp.rf._abc_6362_n7003) );
	NAND2X1 NAND2X1_4796 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7003), .Y(dp.rf._abc_6362_n7004) );
	INVX1 INVX1_164 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<16>), .Y(dp.rf._abc_6362_n7005) );
	NOR2X1 NOR2X1_590 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7005), .Y(dp.rf._abc_6362_n7006) );
	NOR2X1 NOR2X1_591 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7004), .B(dp.rf._abc_6362_n7006), .Y(dp.rf._abc_6362_n7007) );
	OR2X2 OR2X2_52 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7002), .B(dp.rf._abc_6362_n7007), .Y(dp.rf._abc_6362_n7008) );
	NAND2X1 NAND2X1_4797 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7008), .Y(dp.rf._abc_6362_n7009) );
	AND2X2 AND2X2_215 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7009), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7010) );
	NAND2X1 NAND2X1_4798 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6998), .B(dp.rf._abc_6362_n7010), .Y(dp.rf._abc_6362_n7011) );
	NAND2X1 NAND2X1_4799 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7011), .Y(dp.rf._abc_6362_n7012) );
	NOR2X1 NOR2X1_592 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n6988), .B(dp.rf._abc_6362_n7012), .Y(dp.rf._abc_6362_n7013) );
	NAND2X1 NAND2X1_4800 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<16>), .Y(dp.rf._abc_6362_n7014) );
	NAND2X1 NAND2X1_4801 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7014), .Y(dp.rf._abc_6362_n7015) );
	INVX1 INVX1_165 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<16>), .Y(dp.rf._abc_6362_n7016) );
	NOR2X1 NOR2X1_593 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7016), .Y(dp.rf._abc_6362_n7017) );
	NOR2X1 NOR2X1_594 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7015), .B(dp.rf._abc_6362_n7017), .Y(dp.rf._abc_6362_n7018) );
	NAND2X1 NAND2X1_4802 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<16>), .Y(dp.rf._abc_6362_n7019) );
	NAND2X1 NAND2X1_4803 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7019), .Y(dp.rf._abc_6362_n7020) );
	INVX1 INVX1_166 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<16>), .Y(dp.rf._abc_6362_n7021) );
	NOR2X1 NOR2X1_595 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7021), .Y(dp.rf._abc_6362_n7022) );
	NOR2X1 NOR2X1_596 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7020), .B(dp.rf._abc_6362_n7022), .Y(dp.rf._abc_6362_n7023) );
	OR2X2 OR2X2_53 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7018), .B(dp.rf._abc_6362_n7023), .Y(dp.rf._abc_6362_n7024) );
	NAND2X1 NAND2X1_4804 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7024), .Y(dp.rf._abc_6362_n7025) );
	NAND2X1 NAND2X1_4805 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<16>), .Y(dp.rf._abc_6362_n7026) );
	NAND2X1 NAND2X1_4806 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7026), .Y(dp.rf._abc_6362_n7027) );
	INVX1 INVX1_167 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<16>), .Y(dp.rf._abc_6362_n7028) );
	NOR2X1 NOR2X1_597 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7028), .Y(dp.rf._abc_6362_n7029) );
	NOR2X1 NOR2X1_598 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7027), .B(dp.rf._abc_6362_n7029), .Y(dp.rf._abc_6362_n7030) );
	NAND2X1 NAND2X1_4807 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<16>), .Y(dp.rf._abc_6362_n7031) );
	NAND2X1 NAND2X1_4808 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7031), .Y(dp.rf._abc_6362_n7032) );
	INVX1 INVX1_168 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<16>), .Y(dp.rf._abc_6362_n7033) );
	NOR2X1 NOR2X1_599 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7033), .Y(dp.rf._abc_6362_n7034) );
	NOR2X1 NOR2X1_600 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7032), .B(dp.rf._abc_6362_n7034), .Y(dp.rf._abc_6362_n7035) );
	OR2X2 OR2X2_54 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7030), .B(dp.rf._abc_6362_n7035), .Y(dp.rf._abc_6362_n7036) );
	NAND2X1 NAND2X1_4809 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7036), .Y(dp.rf._abc_6362_n7037) );
	AND2X2 AND2X2_216 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7037), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7038) );
	NAND2X1 NAND2X1_4810 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7025), .B(dp.rf._abc_6362_n7038), .Y(dp.rf._abc_6362_n7039) );
	NAND2X1 NAND2X1_4811 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<16>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7040) );
	NAND2X1 NAND2X1_4812 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<16>), .Y(dp.rf._abc_6362_n7041) );
	AND2X2 AND2X2_217 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7041), .B(instr[22]), .Y(dp.rf._abc_6362_n7042) );
	NAND2X1 NAND2X1_4813 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7040), .B(dp.rf._abc_6362_n7042), .Y(dp.rf._abc_6362_n7043) );
	NAND2X1 NAND2X1_4814 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<16>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7044) );
	NAND2X1 NAND2X1_4815 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<16>), .Y(dp.rf._abc_6362_n7045) );
	AND2X2 AND2X2_218 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7045), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7046) );
	NAND2X1 NAND2X1_4816 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7044), .B(dp.rf._abc_6362_n7046), .Y(dp.rf._abc_6362_n7047) );
	NAND2X1 NAND2X1_4817 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7043), .B(dp.rf._abc_6362_n7047), .Y(dp.rf._abc_6362_n7048) );
	AND2X2 AND2X2_219 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7048), .B(instr[23]), .Y(dp.rf._abc_6362_n7049) );
	NAND2X1 NAND2X1_4818 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<16>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7050) );
	NAND2X1 NAND2X1_4819 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<16>), .Y(dp.rf._abc_6362_n7051) );
	AND2X2 AND2X2_220 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7051), .B(instr[22]), .Y(dp.rf._abc_6362_n7052) );
	NAND2X1 NAND2X1_4820 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7050), .B(dp.rf._abc_6362_n7052), .Y(dp.rf._abc_6362_n7053) );
	NAND2X1 NAND2X1_4821 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<16>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7054) );
	NAND2X1 NAND2X1_4822 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<16>), .Y(dp.rf._abc_6362_n7055) );
	AND2X2 AND2X2_221 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7055), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7056) );
	NAND2X1 NAND2X1_4823 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7054), .B(dp.rf._abc_6362_n7056), .Y(dp.rf._abc_6362_n7057) );
	NAND2X1 NAND2X1_4824 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7053), .B(dp.rf._abc_6362_n7057), .Y(dp.rf._abc_6362_n7058) );
	NAND2X1 NAND2X1_4825 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7058), .Y(dp.rf._abc_6362_n7059) );
	NAND2X1 NAND2X1_4826 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7059), .Y(dp.rf._abc_6362_n7060) );
	NOR2X1 NOR2X1_601 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7049), .B(dp.rf._abc_6362_n7060), .Y(dp.rf._abc_6362_n7061) );
	NOR2X1 NOR2X1_602 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7061), .Y(dp.rf._abc_6362_n7062) );
	NAND2X1 NAND2X1_4827 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7039), .B(dp.rf._abc_6362_n7062), .Y(dp.rf._abc_6362_n7063) );
	NAND2X1 NAND2X1_4828 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n7063), .Y(dp.rf._abc_6362_n7064) );
	NOR2X1 NOR2X1_603 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7013), .B(dp.rf._abc_6362_n7064), .Y(dp.srca_16_) );
	NAND2X1 NAND2X1_4829 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<17>), .Y(dp.rf._abc_6362_n7066) );
	NAND2X1 NAND2X1_4830 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<17>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7067) );
	NAND2X1 NAND2X1_4831 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7066), .B(dp.rf._abc_6362_n7067), .Y(dp.rf._abc_6362_n7068) );
	NAND2X1 NAND2X1_4832 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7068), .Y(dp.rf._abc_6362_n7069) );
	NAND2X1 NAND2X1_4833 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<17>), .Y(dp.rf._abc_6362_n7070) );
	NAND2X1 NAND2X1_4834 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<17>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7071) );
	NAND2X1 NAND2X1_4835 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7070), .B(dp.rf._abc_6362_n7071), .Y(dp.rf._abc_6362_n7072) );
	NAND2X1 NAND2X1_4836 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7072), .Y(dp.rf._abc_6362_n7073) );
	NAND2X1 NAND2X1_4837 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7069), .B(dp.rf._abc_6362_n7073), .Y(dp.rf._abc_6362_n7074) );
	NOR2X1 NOR2X1_604 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7074), .Y(dp.rf._abc_6362_n7075) );
	NAND2X1 NAND2X1_4838 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<17>), .Y(dp.rf._abc_6362_n7076) );
	NAND2X1 NAND2X1_4839 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<17>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7077) );
	NAND2X1 NAND2X1_4840 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7076), .B(dp.rf._abc_6362_n7077), .Y(dp.rf._abc_6362_n7078) );
	NAND2X1 NAND2X1_4841 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7078), .Y(dp.rf._abc_6362_n7079) );
	NAND2X1 NAND2X1_4842 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<17>), .Y(dp.rf._abc_6362_n7080) );
	NAND2X1 NAND2X1_4843 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<17>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7081) );
	NAND2X1 NAND2X1_4844 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7080), .B(dp.rf._abc_6362_n7081), .Y(dp.rf._abc_6362_n7082) );
	NAND2X1 NAND2X1_4845 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7082), .Y(dp.rf._abc_6362_n7083) );
	AND2X2 AND2X2_222 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7079), .B(dp.rf._abc_6362_n7083), .Y(dp.rf._abc_6362_n7084) );
	NAND2X1 NAND2X1_4846 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7084), .Y(dp.rf._abc_6362_n7085) );
	NAND2X1 NAND2X1_4847 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n7085), .Y(dp.rf._abc_6362_n7086) );
	NOR2X1 NOR2X1_605 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7075), .B(dp.rf._abc_6362_n7086), .Y(dp.rf._abc_6362_n7087) );
	NAND2X1 NAND2X1_4848 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<17>), .Y(dp.rf._abc_6362_n7088) );
	NAND2X1 NAND2X1_4849 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7088), .Y(dp.rf._abc_6362_n7089) );
	INVX1 INVX1_169 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<17>), .Y(dp.rf._abc_6362_n7090) );
	NOR2X1 NOR2X1_606 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7090), .Y(dp.rf._abc_6362_n7091) );
	NOR2X1 NOR2X1_607 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7089), .B(dp.rf._abc_6362_n7091), .Y(dp.rf._abc_6362_n7092) );
	NAND2X1 NAND2X1_4850 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<17>), .Y(dp.rf._abc_6362_n7093) );
	NAND2X1 NAND2X1_4851 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7093), .Y(dp.rf._abc_6362_n7094) );
	INVX1 INVX1_170 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<17>), .Y(dp.rf._abc_6362_n7095) );
	NOR2X1 NOR2X1_608 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7095), .Y(dp.rf._abc_6362_n7096) );
	NOR2X1 NOR2X1_609 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7094), .B(dp.rf._abc_6362_n7096), .Y(dp.rf._abc_6362_n7097) );
	NOR2X1 NOR2X1_610 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7092), .B(dp.rf._abc_6362_n7097), .Y(dp.rf._abc_6362_n7098) );
	NAND2X1 NAND2X1_4852 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7098), .Y(dp.rf._abc_6362_n7099) );
	NAND2X1 NAND2X1_4853 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<17>), .Y(dp.rf._abc_6362_n7100) );
	NAND2X1 NAND2X1_4854 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7100), .Y(dp.rf._abc_6362_n7101) );
	INVX1 INVX1_171 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<17>), .Y(dp.rf._abc_6362_n7102) );
	NOR2X1 NOR2X1_611 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7102), .Y(dp.rf._abc_6362_n7103) );
	NOR2X1 NOR2X1_612 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7101), .B(dp.rf._abc_6362_n7103), .Y(dp.rf._abc_6362_n7104) );
	NAND2X1 NAND2X1_4855 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<17>), .Y(dp.rf._abc_6362_n7105) );
	NAND2X1 NAND2X1_4856 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7105), .Y(dp.rf._abc_6362_n7106) );
	INVX1 INVX1_172 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<17>), .Y(dp.rf._abc_6362_n7107) );
	NOR2X1 NOR2X1_613 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7107), .Y(dp.rf._abc_6362_n7108) );
	NOR2X1 NOR2X1_614 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7106), .B(dp.rf._abc_6362_n7108), .Y(dp.rf._abc_6362_n7109) );
	NOR2X1 NOR2X1_615 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7104), .B(dp.rf._abc_6362_n7109), .Y(dp.rf._abc_6362_n7110) );
	NAND2X1 NAND2X1_4857 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7110), .Y(dp.rf._abc_6362_n7111) );
	NAND2X1 NAND2X1_4858 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7099), .B(dp.rf._abc_6362_n7111), .Y(dp.rf._abc_6362_n7112) );
	NAND2X1 NAND2X1_4859 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7112), .Y(dp.rf._abc_6362_n7113) );
	NAND2X1 NAND2X1_4860 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7113), .Y(dp.rf._abc_6362_n7114) );
	NOR2X1 NOR2X1_616 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7087), .B(dp.rf._abc_6362_n7114), .Y(dp.rf._abc_6362_n7115) );
	NAND2X1 NAND2X1_4861 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<17>), .Y(dp.rf._abc_6362_n7116) );
	NAND2X1 NAND2X1_4862 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7116), .Y(dp.rf._abc_6362_n7117) );
	INVX1 INVX1_173 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<17>), .Y(dp.rf._abc_6362_n7118) );
	NOR2X1 NOR2X1_617 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7118), .Y(dp.rf._abc_6362_n7119) );
	NOR2X1 NOR2X1_618 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7117), .B(dp.rf._abc_6362_n7119), .Y(dp.rf._abc_6362_n7120) );
	NAND2X1 NAND2X1_4863 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<17>), .Y(dp.rf._abc_6362_n7121) );
	NAND2X1 NAND2X1_4864 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7121), .Y(dp.rf._abc_6362_n7122) );
	INVX1 INVX1_174 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<17>), .Y(dp.rf._abc_6362_n7123) );
	NOR2X1 NOR2X1_619 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7123), .Y(dp.rf._abc_6362_n7124) );
	NOR2X1 NOR2X1_620 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7122), .B(dp.rf._abc_6362_n7124), .Y(dp.rf._abc_6362_n7125) );
	OR2X2 OR2X2_55 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7120), .B(dp.rf._abc_6362_n7125), .Y(dp.rf._abc_6362_n7126) );
	NAND2X1 NAND2X1_4865 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7126), .Y(dp.rf._abc_6362_n7127) );
	NAND2X1 NAND2X1_4866 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<17>), .Y(dp.rf._abc_6362_n7128) );
	NAND2X1 NAND2X1_4867 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7128), .Y(dp.rf._abc_6362_n7129) );
	INVX1 INVX1_175 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<17>), .Y(dp.rf._abc_6362_n7130) );
	NOR2X1 NOR2X1_621 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7130), .Y(dp.rf._abc_6362_n7131) );
	NOR2X1 NOR2X1_622 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7129), .B(dp.rf._abc_6362_n7131), .Y(dp.rf._abc_6362_n7132) );
	NAND2X1 NAND2X1_4868 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<17>), .Y(dp.rf._abc_6362_n7133) );
	NAND2X1 NAND2X1_4869 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7133), .Y(dp.rf._abc_6362_n7134) );
	INVX1 INVX1_176 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<17>), .Y(dp.rf._abc_6362_n7135) );
	NOR2X1 NOR2X1_623 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7135), .Y(dp.rf._abc_6362_n7136) );
	NOR2X1 NOR2X1_624 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7134), .B(dp.rf._abc_6362_n7136), .Y(dp.rf._abc_6362_n7137) );
	OR2X2 OR2X2_56 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7132), .B(dp.rf._abc_6362_n7137), .Y(dp.rf._abc_6362_n7138) );
	NAND2X1 NAND2X1_4870 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7138), .Y(dp.rf._abc_6362_n7139) );
	AND2X2 AND2X2_223 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7139), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7140) );
	NAND2X1 NAND2X1_4871 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7127), .B(dp.rf._abc_6362_n7140), .Y(dp.rf._abc_6362_n7141) );
	NAND2X1 NAND2X1_4872 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<17>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7142) );
	NAND2X1 NAND2X1_4873 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<17>), .Y(dp.rf._abc_6362_n7143) );
	AND2X2 AND2X2_224 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7143), .B(instr[22]), .Y(dp.rf._abc_6362_n7144) );
	NAND2X1 NAND2X1_4874 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7142), .B(dp.rf._abc_6362_n7144), .Y(dp.rf._abc_6362_n7145) );
	NAND2X1 NAND2X1_4875 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<17>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7146) );
	NAND2X1 NAND2X1_4876 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<17>), .Y(dp.rf._abc_6362_n7147) );
	AND2X2 AND2X2_225 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7147), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7148) );
	NAND2X1 NAND2X1_4877 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7146), .B(dp.rf._abc_6362_n7148), .Y(dp.rf._abc_6362_n7149) );
	NAND2X1 NAND2X1_4878 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7145), .B(dp.rf._abc_6362_n7149), .Y(dp.rf._abc_6362_n7150) );
	AND2X2 AND2X2_226 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7150), .B(instr[23]), .Y(dp.rf._abc_6362_n7151) );
	NAND2X1 NAND2X1_4879 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<17>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7152) );
	NAND2X1 NAND2X1_4880 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<17>), .Y(dp.rf._abc_6362_n7153) );
	AND2X2 AND2X2_227 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7153), .B(instr[22]), .Y(dp.rf._abc_6362_n7154) );
	NAND2X1 NAND2X1_4881 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7152), .B(dp.rf._abc_6362_n7154), .Y(dp.rf._abc_6362_n7155) );
	NAND2X1 NAND2X1_4882 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<17>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7156) );
	NAND2X1 NAND2X1_4883 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<17>), .Y(dp.rf._abc_6362_n7157) );
	AND2X2 AND2X2_228 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7157), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7158) );
	NAND2X1 NAND2X1_4884 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7156), .B(dp.rf._abc_6362_n7158), .Y(dp.rf._abc_6362_n7159) );
	NAND2X1 NAND2X1_4885 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7155), .B(dp.rf._abc_6362_n7159), .Y(dp.rf._abc_6362_n7160) );
	NAND2X1 NAND2X1_4886 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7160), .Y(dp.rf._abc_6362_n7161) );
	NAND2X1 NAND2X1_4887 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7161), .Y(dp.rf._abc_6362_n7162) );
	NOR2X1 NOR2X1_625 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7151), .B(dp.rf._abc_6362_n7162), .Y(dp.rf._abc_6362_n7163) );
	NOR2X1 NOR2X1_626 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7163), .Y(dp.rf._abc_6362_n7164) );
	NAND2X1 NAND2X1_4888 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7141), .B(dp.rf._abc_6362_n7164), .Y(dp.rf._abc_6362_n7165) );
	NAND2X1 NAND2X1_4889 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n7165), .Y(dp.rf._abc_6362_n7166) );
	NOR2X1 NOR2X1_627 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7115), .B(dp.rf._abc_6362_n7166), .Y(dp.srca_17_) );
	NAND2X1 NAND2X1_4890 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<18>), .Y(dp.rf._abc_6362_n7168) );
	NAND2X1 NAND2X1_4891 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7168), .Y(dp.rf._abc_6362_n7169) );
	INVX1 INVX1_177 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<18>), .Y(dp.rf._abc_6362_n7170) );
	NOR2X1 NOR2X1_628 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7170), .Y(dp.rf._abc_6362_n7171) );
	NOR2X1 NOR2X1_629 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7169), .B(dp.rf._abc_6362_n7171), .Y(dp.rf._abc_6362_n7172) );
	NAND2X1 NAND2X1_4892 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<18>), .Y(dp.rf._abc_6362_n7173) );
	NAND2X1 NAND2X1_4893 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7173), .Y(dp.rf._abc_6362_n7174) );
	INVX1 INVX1_178 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<18>), .Y(dp.rf._abc_6362_n7175) );
	NOR2X1 NOR2X1_630 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7175), .Y(dp.rf._abc_6362_n7176) );
	NOR2X1 NOR2X1_631 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7174), .B(dp.rf._abc_6362_n7176), .Y(dp.rf._abc_6362_n7177) );
	NOR2X1 NOR2X1_632 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7172), .B(dp.rf._abc_6362_n7177), .Y(dp.rf._abc_6362_n7178) );
	NAND2X1 NAND2X1_4894 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7178), .Y(dp.rf._abc_6362_n7179) );
	NAND2X1 NAND2X1_4895 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<18>), .Y(dp.rf._abc_6362_n7180) );
	NAND2X1 NAND2X1_4896 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7180), .Y(dp.rf._abc_6362_n7181) );
	INVX1 INVX1_179 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<18>), .Y(dp.rf._abc_6362_n7182) );
	NOR2X1 NOR2X1_633 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7182), .Y(dp.rf._abc_6362_n7183) );
	NOR2X1 NOR2X1_634 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7181), .B(dp.rf._abc_6362_n7183), .Y(dp.rf._abc_6362_n7184) );
	NAND2X1 NAND2X1_4897 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<18>), .Y(dp.rf._abc_6362_n7185) );
	NAND2X1 NAND2X1_4898 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7185), .Y(dp.rf._abc_6362_n7186) );
	INVX1 INVX1_180 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<18>), .Y(dp.rf._abc_6362_n7187) );
	NOR2X1 NOR2X1_635 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7187), .Y(dp.rf._abc_6362_n7188) );
	NOR2X1 NOR2X1_636 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7186), .B(dp.rf._abc_6362_n7188), .Y(dp.rf._abc_6362_n7189) );
	NOR2X1 NOR2X1_637 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7184), .B(dp.rf._abc_6362_n7189), .Y(dp.rf._abc_6362_n7190) );
	NAND2X1 NAND2X1_4899 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7190), .Y(dp.rf._abc_6362_n7191) );
	NAND2X1 NAND2X1_4900 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7179), .B(dp.rf._abc_6362_n7191), .Y(dp.rf._abc_6362_n7192) );
	NAND2X1 NAND2X1_4901 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7192), .Y(dp.rf._abc_6362_n7193) );
	NAND2X1 NAND2X1_4902 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<18>), .Y(dp.rf._abc_6362_n7194) );
	NAND2X1 NAND2X1_4903 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<18>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7195) );
	NAND2X1 NAND2X1_4904 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7194), .B(dp.rf._abc_6362_n7195), .Y(dp.rf._abc_6362_n7196) );
	NAND2X1 NAND2X1_4905 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7196), .Y(dp.rf._abc_6362_n7197) );
	NAND2X1 NAND2X1_4906 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<18>), .Y(dp.rf._abc_6362_n7198) );
	NAND2X1 NAND2X1_4907 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<18>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7199) );
	NAND2X1 NAND2X1_4908 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7198), .B(dp.rf._abc_6362_n7199), .Y(dp.rf._abc_6362_n7200) );
	NAND2X1 NAND2X1_4909 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7200), .Y(dp.rf._abc_6362_n7201) );
	AND2X2 AND2X2_229 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7197), .B(dp.rf._abc_6362_n7201), .Y(dp.rf._abc_6362_n7202) );
	NAND2X1 NAND2X1_4910 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7202), .Y(dp.rf._abc_6362_n7203) );
	NAND2X1 NAND2X1_4911 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<18>), .Y(dp.rf._abc_6362_n7204) );
	NAND2X1 NAND2X1_4912 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7204), .Y(dp.rf._abc_6362_n7205) );
	AND2X2 AND2X2_230 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf.rf_2_<18>), .Y(dp.rf._abc_6362_n7206) );
	NOR2X1 NOR2X1_638 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7205), .B(dp.rf._abc_6362_n7206), .Y(dp.rf._abc_6362_n7207) );
	NAND2X1 NAND2X1_4913 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<18>), .Y(dp.rf._abc_6362_n7208) );
	NAND2X1 NAND2X1_4914 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7208), .Y(dp.rf._abc_6362_n7209) );
	INVX1 INVX1_181 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<18>), .Y(dp.rf._abc_6362_n7210) );
	NOR2X1 NOR2X1_639 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7210), .Y(dp.rf._abc_6362_n7211) );
	NOR2X1 NOR2X1_640 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7209), .B(dp.rf._abc_6362_n7211), .Y(dp.rf._abc_6362_n7212) );
	OR2X2 OR2X2_57 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7207), .B(dp.rf._abc_6362_n7212), .Y(dp.rf._abc_6362_n7213) );
	NAND2X1 NAND2X1_4915 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7213), .Y(dp.rf._abc_6362_n7214) );
	AND2X2 AND2X2_231 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7214), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7215) );
	NAND2X1 NAND2X1_4916 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7203), .B(dp.rf._abc_6362_n7215), .Y(dp.rf._abc_6362_n7216) );
	NAND2X1 NAND2X1_4917 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7193), .B(dp.rf._abc_6362_n7216), .Y(dp.rf._abc_6362_n7217) );
	NOR2X1 NOR2X1_641 ( .gnd(gnd), .vdd(vdd), .A(instr[25]), .B(dp.rf._abc_6362_n7217), .Y(dp.rf._abc_6362_n7218) );
	NAND2X1 NAND2X1_4918 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<18>), .Y(dp.rf._abc_6362_n7219) );
	NAND2X1 NAND2X1_4919 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7219), .Y(dp.rf._abc_6362_n7220) );
	INVX1 INVX1_182 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<18>), .Y(dp.rf._abc_6362_n7221) );
	NOR2X1 NOR2X1_642 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7221), .Y(dp.rf._abc_6362_n7222) );
	NOR2X1 NOR2X1_643 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7220), .B(dp.rf._abc_6362_n7222), .Y(dp.rf._abc_6362_n7223) );
	NAND2X1 NAND2X1_4920 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<18>), .Y(dp.rf._abc_6362_n7224) );
	NAND2X1 NAND2X1_4921 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7224), .Y(dp.rf._abc_6362_n7225) );
	INVX1 INVX1_183 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<18>), .Y(dp.rf._abc_6362_n7226) );
	NOR2X1 NOR2X1_644 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7226), .Y(dp.rf._abc_6362_n7227) );
	NOR2X1 NOR2X1_645 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7225), .B(dp.rf._abc_6362_n7227), .Y(dp.rf._abc_6362_n7228) );
	OR2X2 OR2X2_58 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7223), .B(dp.rf._abc_6362_n7228), .Y(dp.rf._abc_6362_n7229) );
	NAND2X1 NAND2X1_4922 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7229), .Y(dp.rf._abc_6362_n7230) );
	NAND2X1 NAND2X1_4923 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<18>), .Y(dp.rf._abc_6362_n7231) );
	NAND2X1 NAND2X1_4924 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7231), .Y(dp.rf._abc_6362_n7232) );
	INVX1 INVX1_184 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<18>), .Y(dp.rf._abc_6362_n7233) );
	NOR2X1 NOR2X1_646 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7233), .Y(dp.rf._abc_6362_n7234) );
	NOR2X1 NOR2X1_647 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7232), .B(dp.rf._abc_6362_n7234), .Y(dp.rf._abc_6362_n7235) );
	NAND2X1 NAND2X1_4925 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<18>), .Y(dp.rf._abc_6362_n7236) );
	NAND2X1 NAND2X1_4926 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7236), .Y(dp.rf._abc_6362_n7237) );
	INVX1 INVX1_185 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<18>), .Y(dp.rf._abc_6362_n7238) );
	NOR2X1 NOR2X1_648 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7238), .Y(dp.rf._abc_6362_n7239) );
	NOR2X1 NOR2X1_649 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7237), .B(dp.rf._abc_6362_n7239), .Y(dp.rf._abc_6362_n7240) );
	OR2X2 OR2X2_59 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7235), .B(dp.rf._abc_6362_n7240), .Y(dp.rf._abc_6362_n7241) );
	NAND2X1 NAND2X1_4927 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7241), .Y(dp.rf._abc_6362_n7242) );
	AND2X2 AND2X2_232 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7242), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7243) );
	NAND2X1 NAND2X1_4928 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7230), .B(dp.rf._abc_6362_n7243), .Y(dp.rf._abc_6362_n7244) );
	NAND2X1 NAND2X1_4929 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<18>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7245) );
	NAND2X1 NAND2X1_4930 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<18>), .Y(dp.rf._abc_6362_n7246) );
	AND2X2 AND2X2_233 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7246), .B(instr[22]), .Y(dp.rf._abc_6362_n7247) );
	NAND2X1 NAND2X1_4931 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7245), .B(dp.rf._abc_6362_n7247), .Y(dp.rf._abc_6362_n7248) );
	NAND2X1 NAND2X1_4932 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<18>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7249) );
	NAND2X1 NAND2X1_4933 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<18>), .Y(dp.rf._abc_6362_n7250) );
	AND2X2 AND2X2_234 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7250), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7251) );
	NAND2X1 NAND2X1_4934 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7249), .B(dp.rf._abc_6362_n7251), .Y(dp.rf._abc_6362_n7252) );
	NAND2X1 NAND2X1_4935 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7248), .B(dp.rf._abc_6362_n7252), .Y(dp.rf._abc_6362_n7253) );
	AND2X2 AND2X2_235 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7253), .B(instr[23]), .Y(dp.rf._abc_6362_n7254) );
	NAND2X1 NAND2X1_4936 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<18>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7255) );
	NAND2X1 NAND2X1_4937 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<18>), .Y(dp.rf._abc_6362_n7256) );
	AND2X2 AND2X2_236 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7256), .B(instr[22]), .Y(dp.rf._abc_6362_n7257) );
	NAND2X1 NAND2X1_4938 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7255), .B(dp.rf._abc_6362_n7257), .Y(dp.rf._abc_6362_n7258) );
	NAND2X1 NAND2X1_4939 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<18>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7259) );
	NAND2X1 NAND2X1_4940 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<18>), .Y(dp.rf._abc_6362_n7260) );
	AND2X2 AND2X2_237 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7260), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7261) );
	NAND2X1 NAND2X1_4941 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7259), .B(dp.rf._abc_6362_n7261), .Y(dp.rf._abc_6362_n7262) );
	NAND2X1 NAND2X1_4942 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7258), .B(dp.rf._abc_6362_n7262), .Y(dp.rf._abc_6362_n7263) );
	NAND2X1 NAND2X1_4943 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7263), .Y(dp.rf._abc_6362_n7264) );
	NAND2X1 NAND2X1_4944 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7264), .Y(dp.rf._abc_6362_n7265) );
	NOR2X1 NOR2X1_650 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7254), .B(dp.rf._abc_6362_n7265), .Y(dp.rf._abc_6362_n7266) );
	NOR2X1 NOR2X1_651 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7266), .Y(dp.rf._abc_6362_n7267) );
	NAND2X1 NAND2X1_4945 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7244), .B(dp.rf._abc_6362_n7267), .Y(dp.rf._abc_6362_n7268) );
	NAND2X1 NAND2X1_4946 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n7268), .Y(dp.rf._abc_6362_n7269) );
	NOR2X1 NOR2X1_652 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7218), .B(dp.rf._abc_6362_n7269), .Y(dp.srca_18_) );
	NAND2X1 NAND2X1_4947 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<19>), .Y(dp.rf._abc_6362_n7271) );
	NAND2X1 NAND2X1_4948 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7272) );
	NAND2X1 NAND2X1_4949 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7271), .B(dp.rf._abc_6362_n7272), .Y(dp.rf._abc_6362_n7273) );
	NAND2X1 NAND2X1_4950 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7273), .Y(dp.rf._abc_6362_n7274) );
	NAND2X1 NAND2X1_4951 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<19>), .Y(dp.rf._abc_6362_n7275) );
	NAND2X1 NAND2X1_4952 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7276) );
	NAND2X1 NAND2X1_4953 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7275), .B(dp.rf._abc_6362_n7276), .Y(dp.rf._abc_6362_n7277) );
	NAND2X1 NAND2X1_4954 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7277), .Y(dp.rf._abc_6362_n7278) );
	NAND2X1 NAND2X1_4955 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7274), .B(dp.rf._abc_6362_n7278), .Y(dp.rf._abc_6362_n7279) );
	NOR2X1 NOR2X1_653 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7279), .Y(dp.rf._abc_6362_n7280) );
	NAND2X1 NAND2X1_4956 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<19>), .Y(dp.rf._abc_6362_n7281) );
	NAND2X1 NAND2X1_4957 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7282) );
	NAND2X1 NAND2X1_4958 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7281), .B(dp.rf._abc_6362_n7282), .Y(dp.rf._abc_6362_n7283) );
	NAND2X1 NAND2X1_4959 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7283), .Y(dp.rf._abc_6362_n7284) );
	NAND2X1 NAND2X1_4960 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<19>), .Y(dp.rf._abc_6362_n7285) );
	NAND2X1 NAND2X1_4961 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7286) );
	NAND2X1 NAND2X1_4962 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7285), .B(dp.rf._abc_6362_n7286), .Y(dp.rf._abc_6362_n7287) );
	NAND2X1 NAND2X1_4963 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7287), .Y(dp.rf._abc_6362_n7288) );
	AND2X2 AND2X2_238 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7284), .B(dp.rf._abc_6362_n7288), .Y(dp.rf._abc_6362_n7289) );
	NAND2X1 NAND2X1_4964 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7289), .Y(dp.rf._abc_6362_n7290) );
	NAND2X1 NAND2X1_4965 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n7290), .Y(dp.rf._abc_6362_n7291) );
	NOR2X1 NOR2X1_654 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7280), .B(dp.rf._abc_6362_n7291), .Y(dp.rf._abc_6362_n7292) );
	NAND2X1 NAND2X1_4966 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<19>), .Y(dp.rf._abc_6362_n7293) );
	NAND2X1 NAND2X1_4967 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7294) );
	NAND2X1 NAND2X1_4968 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7293), .B(dp.rf._abc_6362_n7294), .Y(dp.rf._abc_6362_n7295) );
	NAND2X1 NAND2X1_4969 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7295), .Y(dp.rf._abc_6362_n7296) );
	NAND2X1 NAND2X1_4970 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<19>), .Y(dp.rf._abc_6362_n7297) );
	NAND2X1 NAND2X1_4971 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7298) );
	NAND2X1 NAND2X1_4972 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7297), .B(dp.rf._abc_6362_n7298), .Y(dp.rf._abc_6362_n7299) );
	NAND2X1 NAND2X1_4973 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7299), .Y(dp.rf._abc_6362_n7300) );
	AND2X2 AND2X2_239 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7296), .B(dp.rf._abc_6362_n7300), .Y(dp.rf._abc_6362_n7301) );
	NAND2X1 NAND2X1_4974 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7301), .Y(dp.rf._abc_6362_n7302) );
	NAND2X1 NAND2X1_4975 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<19>), .Y(dp.rf._abc_6362_n7303) );
	NAND2X1 NAND2X1_4976 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7303), .Y(dp.rf._abc_6362_n7304) );
	AND2X2 AND2X2_240 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf.rf_10_<19>), .Y(dp.rf._abc_6362_n7305) );
	NOR2X1 NOR2X1_655 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7304), .B(dp.rf._abc_6362_n7305), .Y(dp.rf._abc_6362_n7306) );
	NAND2X1 NAND2X1_4977 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<19>), .Y(dp.rf._abc_6362_n7307) );
	NAND2X1 NAND2X1_4978 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7307), .Y(dp.rf._abc_6362_n7308) );
	INVX1 INVX1_186 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<19>), .Y(dp.rf._abc_6362_n7309) );
	NOR2X1 NOR2X1_656 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7309), .Y(dp.rf._abc_6362_n7310) );
	NOR2X1 NOR2X1_657 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7308), .B(dp.rf._abc_6362_n7310), .Y(dp.rf._abc_6362_n7311) );
	OR2X2 OR2X2_60 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7306), .B(dp.rf._abc_6362_n7311), .Y(dp.rf._abc_6362_n7312) );
	NAND2X1 NAND2X1_4979 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7312), .Y(dp.rf._abc_6362_n7313) );
	AND2X2 AND2X2_241 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7313), .B(instr[24]), .Y(dp.rf._abc_6362_n7314) );
	NAND2X1 NAND2X1_4980 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7302), .B(dp.rf._abc_6362_n7314), .Y(dp.rf._abc_6362_n7315) );
	NAND2X1 NAND2X1_4981 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7315), .Y(dp.rf._abc_6362_n7316) );
	NOR2X1 NOR2X1_658 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7292), .B(dp.rf._abc_6362_n7316), .Y(dp.rf._abc_6362_n7317) );
	NAND2X1 NAND2X1_4982 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<19>), .Y(dp.rf._abc_6362_n7318) );
	NAND2X1 NAND2X1_4983 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7319) );
	NAND2X1 NAND2X1_4984 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7318), .B(dp.rf._abc_6362_n7319), .Y(dp.rf._abc_6362_n7320) );
	NAND2X1 NAND2X1_4985 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7320), .Y(dp.rf._abc_6362_n7321) );
	NAND2X1 NAND2X1_4986 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<19>), .Y(dp.rf._abc_6362_n7322) );
	NAND2X1 NAND2X1_4987 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7323) );
	NAND2X1 NAND2X1_4988 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7322), .B(dp.rf._abc_6362_n7323), .Y(dp.rf._abc_6362_n7324) );
	NAND2X1 NAND2X1_4989 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7324), .Y(dp.rf._abc_6362_n7325) );
	AND2X2 AND2X2_242 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7321), .B(dp.rf._abc_6362_n7325), .Y(dp.rf._abc_6362_n7326) );
	NAND2X1 NAND2X1_4990 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7326), .Y(dp.rf._abc_6362_n7327) );
	NAND2X1 NAND2X1_4991 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<19>), .Y(dp.rf._abc_6362_n7328) );
	NAND2X1 NAND2X1_4992 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7329) );
	NAND2X1 NAND2X1_4993 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7328), .B(dp.rf._abc_6362_n7329), .Y(dp.rf._abc_6362_n7330) );
	NAND2X1 NAND2X1_4994 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7330), .Y(dp.rf._abc_6362_n7331) );
	NAND2X1 NAND2X1_4995 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<19>), .Y(dp.rf._abc_6362_n7332) );
	NAND2X1 NAND2X1_4996 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7333) );
	NAND2X1 NAND2X1_4997 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7332), .B(dp.rf._abc_6362_n7333), .Y(dp.rf._abc_6362_n7334) );
	NAND2X1 NAND2X1_4998 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7334), .Y(dp.rf._abc_6362_n7335) );
	AND2X2 AND2X2_243 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7331), .B(dp.rf._abc_6362_n7335), .Y(dp.rf._abc_6362_n7336) );
	NAND2X1 NAND2X1_4999 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7336), .Y(dp.rf._abc_6362_n7337) );
	AND2X2 AND2X2_244 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7337), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7338) );
	NAND2X1 NAND2X1_5000 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7327), .B(dp.rf._abc_6362_n7338), .Y(dp.rf._abc_6362_n7339) );
	NAND2X1 NAND2X1_5001 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7340) );
	NAND2X1 NAND2X1_5002 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<19>), .Y(dp.rf._abc_6362_n7341) );
	AND2X2 AND2X2_245 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7341), .B(instr[22]), .Y(dp.rf._abc_6362_n7342) );
	NAND2X1 NAND2X1_5003 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7340), .B(dp.rf._abc_6362_n7342), .Y(dp.rf._abc_6362_n7343) );
	NAND2X1 NAND2X1_5004 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7344) );
	NAND2X1 NAND2X1_5005 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<19>), .Y(dp.rf._abc_6362_n7345) );
	AND2X2 AND2X2_246 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7345), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7346) );
	NAND2X1 NAND2X1_5006 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7344), .B(dp.rf._abc_6362_n7346), .Y(dp.rf._abc_6362_n7347) );
	NAND2X1 NAND2X1_5007 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7343), .B(dp.rf._abc_6362_n7347), .Y(dp.rf._abc_6362_n7348) );
	AND2X2 AND2X2_247 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7348), .B(instr[23]), .Y(dp.rf._abc_6362_n7349) );
	NAND2X1 NAND2X1_5008 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7350) );
	NAND2X1 NAND2X1_5009 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<19>), .Y(dp.rf._abc_6362_n7351) );
	AND2X2 AND2X2_248 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7351), .B(instr[22]), .Y(dp.rf._abc_6362_n7352) );
	NAND2X1 NAND2X1_5010 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7350), .B(dp.rf._abc_6362_n7352), .Y(dp.rf._abc_6362_n7353) );
	NAND2X1 NAND2X1_5011 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<19>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7354) );
	NAND2X1 NAND2X1_5012 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<19>), .Y(dp.rf._abc_6362_n7355) );
	AND2X2 AND2X2_249 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7355), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7356) );
	NAND2X1 NAND2X1_5013 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7354), .B(dp.rf._abc_6362_n7356), .Y(dp.rf._abc_6362_n7357) );
	NAND2X1 NAND2X1_5014 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7353), .B(dp.rf._abc_6362_n7357), .Y(dp.rf._abc_6362_n7358) );
	NAND2X1 NAND2X1_5015 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7358), .Y(dp.rf._abc_6362_n7359) );
	NAND2X1 NAND2X1_5016 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7359), .Y(dp.rf._abc_6362_n7360) );
	NOR2X1 NOR2X1_659 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7349), .B(dp.rf._abc_6362_n7360), .Y(dp.rf._abc_6362_n7361) );
	NOR2X1 NOR2X1_660 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7361), .Y(dp.rf._abc_6362_n7362) );
	NAND2X1 NAND2X1_5017 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7339), .B(dp.rf._abc_6362_n7362), .Y(dp.rf._abc_6362_n7363) );
	NAND2X1 NAND2X1_5018 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n7363), .Y(dp.rf._abc_6362_n7364) );
	NOR2X1 NOR2X1_661 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7317), .B(dp.rf._abc_6362_n7364), .Y(dp.srca_19_) );
	NAND2X1 NAND2X1_5019 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<20>), .Y(dp.rf._abc_6362_n7366) );
	NAND2X1 NAND2X1_5020 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7367) );
	NAND2X1 NAND2X1_5021 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7366), .B(dp.rf._abc_6362_n7367), .Y(dp.rf._abc_6362_n7368) );
	NAND2X1 NAND2X1_5022 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7368), .Y(dp.rf._abc_6362_n7369) );
	NAND2X1 NAND2X1_5023 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<20>), .Y(dp.rf._abc_6362_n7370) );
	NAND2X1 NAND2X1_5024 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7371) );
	NAND2X1 NAND2X1_5025 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7370), .B(dp.rf._abc_6362_n7371), .Y(dp.rf._abc_6362_n7372) );
	NAND2X1 NAND2X1_5026 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7372), .Y(dp.rf._abc_6362_n7373) );
	NAND2X1 NAND2X1_5027 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7369), .B(dp.rf._abc_6362_n7373), .Y(dp.rf._abc_6362_n7374) );
	NAND2X1 NAND2X1_5028 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7374), .Y(dp.rf._abc_6362_n7375) );
	NAND2X1 NAND2X1_5029 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<20>), .Y(dp.rf._abc_6362_n7376) );
	NAND2X1 NAND2X1_5030 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7377) );
	NAND2X1 NAND2X1_5031 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7376), .B(dp.rf._abc_6362_n7377), .Y(dp.rf._abc_6362_n7378) );
	NAND2X1 NAND2X1_5032 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7378), .Y(dp.rf._abc_6362_n7379) );
	NAND2X1 NAND2X1_5033 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<20>), .Y(dp.rf._abc_6362_n7380) );
	NAND2X1 NAND2X1_5034 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7381) );
	NAND2X1 NAND2X1_5035 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7380), .B(dp.rf._abc_6362_n7381), .Y(dp.rf._abc_6362_n7382) );
	NAND2X1 NAND2X1_5036 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7382), .Y(dp.rf._abc_6362_n7383) );
	NAND2X1 NAND2X1_5037 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7379), .B(dp.rf._abc_6362_n7383), .Y(dp.rf._abc_6362_n7384) );
	NAND2X1 NAND2X1_5038 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7384), .Y(dp.rf._abc_6362_n7385) );
	NAND2X1 NAND2X1_5039 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7375), .B(dp.rf._abc_6362_n7385), .Y(dp.rf._abc_6362_n7386) );
	NAND2X1 NAND2X1_5040 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7386), .Y(dp.rf._abc_6362_n7387) );
	NAND2X1 NAND2X1_5041 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<20>), .Y(dp.rf._abc_6362_n7388) );
	NAND2X1 NAND2X1_5042 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7388), .Y(dp.rf._abc_6362_n7389) );
	INVX1 INVX1_187 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<20>), .Y(dp.rf._abc_6362_n7390) );
	NOR2X1 NOR2X1_662 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7390), .Y(dp.rf._abc_6362_n7391) );
	NOR2X1 NOR2X1_663 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7389), .B(dp.rf._abc_6362_n7391), .Y(dp.rf._abc_6362_n7392) );
	NAND2X1 NAND2X1_5043 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<20>), .Y(dp.rf._abc_6362_n7393) );
	NAND2X1 NAND2X1_5044 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7393), .Y(dp.rf._abc_6362_n7394) );
	INVX1 INVX1_188 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<20>), .Y(dp.rf._abc_6362_n7395) );
	NOR2X1 NOR2X1_664 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7395), .Y(dp.rf._abc_6362_n7396) );
	NOR2X1 NOR2X1_665 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7394), .B(dp.rf._abc_6362_n7396), .Y(dp.rf._abc_6362_n7397) );
	OR2X2 OR2X2_61 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7392), .B(dp.rf._abc_6362_n7397), .Y(dp.rf._abc_6362_n7398) );
	NAND2X1 NAND2X1_5045 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7398), .Y(dp.rf._abc_6362_n7399) );
	NAND2X1 NAND2X1_5046 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<20>), .Y(dp.rf._abc_6362_n7400) );
	NAND2X1 NAND2X1_5047 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7400), .Y(dp.rf._abc_6362_n7401) );
	INVX1 INVX1_189 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<20>), .Y(dp.rf._abc_6362_n7402) );
	NOR2X1 NOR2X1_666 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7402), .Y(dp.rf._abc_6362_n7403) );
	NOR2X1 NOR2X1_667 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7401), .B(dp.rf._abc_6362_n7403), .Y(dp.rf._abc_6362_n7404) );
	NAND2X1 NAND2X1_5048 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<20>), .Y(dp.rf._abc_6362_n7405) );
	NAND2X1 NAND2X1_5049 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7405), .Y(dp.rf._abc_6362_n7406) );
	INVX1 INVX1_190 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<20>), .Y(dp.rf._abc_6362_n7407) );
	NOR2X1 NOR2X1_668 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7407), .Y(dp.rf._abc_6362_n7408) );
	NOR2X1 NOR2X1_669 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7406), .B(dp.rf._abc_6362_n7408), .Y(dp.rf._abc_6362_n7409) );
	OR2X2 OR2X2_62 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7404), .B(dp.rf._abc_6362_n7409), .Y(dp.rf._abc_6362_n7410) );
	NAND2X1 NAND2X1_5050 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7410), .Y(dp.rf._abc_6362_n7411) );
	AND2X2 AND2X2_250 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7411), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7412) );
	NAND2X1 NAND2X1_5051 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7399), .B(dp.rf._abc_6362_n7412), .Y(dp.rf._abc_6362_n7413) );
	NAND2X1 NAND2X1_5052 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7387), .B(dp.rf._abc_6362_n7413), .Y(dp.rf._abc_6362_n7414) );
	NOR2X1 NOR2X1_670 ( .gnd(gnd), .vdd(vdd), .A(instr[25]), .B(dp.rf._abc_6362_n7414), .Y(dp.rf._abc_6362_n7415) );
	NAND2X1 NAND2X1_5053 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<20>), .Y(dp.rf._abc_6362_n7416) );
	NAND2X1 NAND2X1_5054 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7417) );
	NAND2X1 NAND2X1_5055 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7416), .B(dp.rf._abc_6362_n7417), .Y(dp.rf._abc_6362_n7418) );
	NAND2X1 NAND2X1_5056 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7418), .Y(dp.rf._abc_6362_n7419) );
	NAND2X1 NAND2X1_5057 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<20>), .Y(dp.rf._abc_6362_n7420) );
	NAND2X1 NAND2X1_5058 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7421) );
	NAND2X1 NAND2X1_5059 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7420), .B(dp.rf._abc_6362_n7421), .Y(dp.rf._abc_6362_n7422) );
	NAND2X1 NAND2X1_5060 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7422), .Y(dp.rf._abc_6362_n7423) );
	NAND2X1 NAND2X1_5061 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7419), .B(dp.rf._abc_6362_n7423), .Y(dp.rf._abc_6362_n7424) );
	NAND2X1 NAND2X1_5062 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7424), .Y(dp.rf._abc_6362_n7425) );
	NAND2X1 NAND2X1_5063 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<20>), .Y(dp.rf._abc_6362_n7426) );
	NAND2X1 NAND2X1_5064 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7427) );
	NAND2X1 NAND2X1_5065 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7426), .B(dp.rf._abc_6362_n7427), .Y(dp.rf._abc_6362_n7428) );
	NAND2X1 NAND2X1_5066 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7428), .Y(dp.rf._abc_6362_n7429) );
	NAND2X1 NAND2X1_5067 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<20>), .Y(dp.rf._abc_6362_n7430) );
	NAND2X1 NAND2X1_5068 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7431) );
	NAND2X1 NAND2X1_5069 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7430), .B(dp.rf._abc_6362_n7431), .Y(dp.rf._abc_6362_n7432) );
	NAND2X1 NAND2X1_5070 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7432), .Y(dp.rf._abc_6362_n7433) );
	NAND2X1 NAND2X1_5071 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7429), .B(dp.rf._abc_6362_n7433), .Y(dp.rf._abc_6362_n7434) );
	NAND2X1 NAND2X1_5072 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7434), .Y(dp.rf._abc_6362_n7435) );
	NAND2X1 NAND2X1_5073 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7425), .B(dp.rf._abc_6362_n7435), .Y(dp.rf._abc_6362_n7436) );
	NAND2X1 NAND2X1_5074 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7436), .Y(dp.rf._abc_6362_n7437) );
	NAND2X1 NAND2X1_5075 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7438) );
	NAND2X1 NAND2X1_5076 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<20>), .Y(dp.rf._abc_6362_n7439) );
	AND2X2 AND2X2_251 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7439), .B(instr[22]), .Y(dp.rf._abc_6362_n7440) );
	NAND2X1 NAND2X1_5077 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7438), .B(dp.rf._abc_6362_n7440), .Y(dp.rf._abc_6362_n7441) );
	NAND2X1 NAND2X1_5078 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7442) );
	NAND2X1 NAND2X1_5079 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<20>), .Y(dp.rf._abc_6362_n7443) );
	AND2X2 AND2X2_252 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7443), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7444) );
	NAND2X1 NAND2X1_5080 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7442), .B(dp.rf._abc_6362_n7444), .Y(dp.rf._abc_6362_n7445) );
	NAND2X1 NAND2X1_5081 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7441), .B(dp.rf._abc_6362_n7445), .Y(dp.rf._abc_6362_n7446) );
	AND2X2 AND2X2_253 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7446), .B(instr[23]), .Y(dp.rf._abc_6362_n7447) );
	NAND2X1 NAND2X1_5082 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7448) );
	NAND2X1 NAND2X1_5083 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<20>), .Y(dp.rf._abc_6362_n7449) );
	AND2X2 AND2X2_254 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7449), .B(instr[22]), .Y(dp.rf._abc_6362_n7450) );
	NAND2X1 NAND2X1_5084 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7448), .B(dp.rf._abc_6362_n7450), .Y(dp.rf._abc_6362_n7451) );
	NAND2X1 NAND2X1_5085 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<20>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7452) );
	NAND2X1 NAND2X1_5086 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<20>), .Y(dp.rf._abc_6362_n7453) );
	AND2X2 AND2X2_255 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7453), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7454) );
	NAND2X1 NAND2X1_5087 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7452), .B(dp.rf._abc_6362_n7454), .Y(dp.rf._abc_6362_n7455) );
	NAND2X1 NAND2X1_5088 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7451), .B(dp.rf._abc_6362_n7455), .Y(dp.rf._abc_6362_n7456) );
	NAND2X1 NAND2X1_5089 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7456), .Y(dp.rf._abc_6362_n7457) );
	NAND2X1 NAND2X1_5090 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n7457), .Y(dp.rf._abc_6362_n7458) );
	NOR2X1 NOR2X1_671 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7447), .B(dp.rf._abc_6362_n7458), .Y(dp.rf._abc_6362_n7459) );
	NOR2X1 NOR2X1_672 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7459), .Y(dp.rf._abc_6362_n7460) );
	NAND2X1 NAND2X1_5091 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7437), .B(dp.rf._abc_6362_n7460), .Y(dp.rf._abc_6362_n7461) );
	NAND2X1 NAND2X1_5092 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n7461), .Y(dp.rf._abc_6362_n7462) );
	NOR2X1 NOR2X1_673 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7415), .B(dp.rf._abc_6362_n7462), .Y(dp.srca_20_) );
	NAND2X1 NAND2X1_5093 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<21>), .Y(dp.rf._abc_6362_n7464) );
	NAND2X1 NAND2X1_5094 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<21>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7465) );
	NAND2X1 NAND2X1_5095 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7464), .B(dp.rf._abc_6362_n7465), .Y(dp.rf._abc_6362_n7466) );
	NAND2X1 NAND2X1_5096 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7466), .Y(dp.rf._abc_6362_n7467) );
	NAND2X1 NAND2X1_5097 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<21>), .Y(dp.rf._abc_6362_n7468) );
	NAND2X1 NAND2X1_5098 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<21>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7469) );
	NAND2X1 NAND2X1_5099 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7468), .B(dp.rf._abc_6362_n7469), .Y(dp.rf._abc_6362_n7470) );
	NAND2X1 NAND2X1_5100 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7470), .Y(dp.rf._abc_6362_n7471) );
	NAND2X1 NAND2X1_5101 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7467), .B(dp.rf._abc_6362_n7471), .Y(dp.rf._abc_6362_n7472) );
	NOR2X1 NOR2X1_674 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7472), .Y(dp.rf._abc_6362_n7473) );
	NAND2X1 NAND2X1_5102 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<21>), .Y(dp.rf._abc_6362_n7474) );
	NAND2X1 NAND2X1_5103 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<21>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7475) );
	NAND2X1 NAND2X1_5104 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7474), .B(dp.rf._abc_6362_n7475), .Y(dp.rf._abc_6362_n7476) );
	NAND2X1 NAND2X1_5105 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7476), .Y(dp.rf._abc_6362_n7477) );
	NAND2X1 NAND2X1_5106 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<21>), .Y(dp.rf._abc_6362_n7478) );
	NAND2X1 NAND2X1_5107 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<21>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7479) );
	NAND2X1 NAND2X1_5108 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7478), .B(dp.rf._abc_6362_n7479), .Y(dp.rf._abc_6362_n7480) );
	NAND2X1 NAND2X1_5109 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7480), .Y(dp.rf._abc_6362_n7481) );
	AND2X2 AND2X2_256 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7477), .B(dp.rf._abc_6362_n7481), .Y(dp.rf._abc_6362_n7482) );
	NAND2X1 NAND2X1_5110 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7482), .Y(dp.rf._abc_6362_n7483) );
	NAND2X1 NAND2X1_5111 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7483), .Y(dp.rf._abc_6362_n7484) );
	NOR2X1 NOR2X1_675 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7473), .B(dp.rf._abc_6362_n7484), .Y(dp.rf._abc_6362_n7485) );
	NAND2X1 NAND2X1_5112 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<21>), .Y(dp.rf._abc_6362_n7486) );
	NAND2X1 NAND2X1_5113 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<21>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7487) );
	NAND2X1 NAND2X1_5114 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7486), .B(dp.rf._abc_6362_n7487), .Y(dp.rf._abc_6362_n7488) );
	NAND2X1 NAND2X1_5115 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7488), .Y(dp.rf._abc_6362_n7489) );
	NAND2X1 NAND2X1_5116 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<21>), .Y(dp.rf._abc_6362_n7490) );
	NAND2X1 NAND2X1_5117 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<21>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7491) );
	NAND2X1 NAND2X1_5118 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7490), .B(dp.rf._abc_6362_n7491), .Y(dp.rf._abc_6362_n7492) );
	NAND2X1 NAND2X1_5119 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7492), .Y(dp.rf._abc_6362_n7493) );
	AND2X2 AND2X2_257 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7489), .B(dp.rf._abc_6362_n7493), .Y(dp.rf._abc_6362_n7494) );
	NAND2X1 NAND2X1_5120 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7494), .Y(dp.rf._abc_6362_n7495) );
	NAND2X1 NAND2X1_5121 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<21>), .Y(dp.rf._abc_6362_n7496) );
	NAND2X1 NAND2X1_5122 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7496), .Y(dp.rf._abc_6362_n7497) );
	AND2X2 AND2X2_258 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf.rf_2_<21>), .Y(dp.rf._abc_6362_n7498) );
	NOR2X1 NOR2X1_676 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7497), .B(dp.rf._abc_6362_n7498), .Y(dp.rf._abc_6362_n7499) );
	NAND2X1 NAND2X1_5123 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<21>), .Y(dp.rf._abc_6362_n7500) );
	NAND2X1 NAND2X1_5124 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7500), .Y(dp.rf._abc_6362_n7501) );
	INVX1 INVX1_191 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<21>), .Y(dp.rf._abc_6362_n7502) );
	NOR2X1 NOR2X1_677 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7502), .Y(dp.rf._abc_6362_n7503) );
	NOR2X1 NOR2X1_678 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7501), .B(dp.rf._abc_6362_n7503), .Y(dp.rf._abc_6362_n7504) );
	OR2X2 OR2X2_63 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7499), .B(dp.rf._abc_6362_n7504), .Y(dp.rf._abc_6362_n7505) );
	NAND2X1 NAND2X1_5125 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7505), .Y(dp.rf._abc_6362_n7506) );
	AND2X2 AND2X2_259 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7506), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7507) );
	NAND2X1 NAND2X1_5126 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7495), .B(dp.rf._abc_6362_n7507), .Y(dp.rf._abc_6362_n7508) );
	NAND2X1 NAND2X1_5127 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7508), .Y(dp.rf._abc_6362_n7509) );
	NOR2X1 NOR2X1_679 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7485), .B(dp.rf._abc_6362_n7509), .Y(dp.rf._abc_6362_n7510) );
	NAND2X1 NAND2X1_5128 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<21>), .Y(dp.rf._abc_6362_n7511) );
	NAND2X1 NAND2X1_5129 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7511), .Y(dp.rf._abc_6362_n7512) );
	INVX1 INVX1_192 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<21>), .Y(dp.rf._abc_6362_n7513) );
	NOR2X1 NOR2X1_680 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7513), .Y(dp.rf._abc_6362_n7514) );
	NOR2X1 NOR2X1_681 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7512), .B(dp.rf._abc_6362_n7514), .Y(dp.rf._abc_6362_n7515) );
	NAND2X1 NAND2X1_5130 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<21>), .Y(dp.rf._abc_6362_n7516) );
	NAND2X1 NAND2X1_5131 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7516), .Y(dp.rf._abc_6362_n7517) );
	INVX1 INVX1_193 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<21>), .Y(dp.rf._abc_6362_n7518) );
	NOR2X1 NOR2X1_682 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7518), .Y(dp.rf._abc_6362_n7519) );
	NOR2X1 NOR2X1_683 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7517), .B(dp.rf._abc_6362_n7519), .Y(dp.rf._abc_6362_n7520) );
	OR2X2 OR2X2_64 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7515), .B(dp.rf._abc_6362_n7520), .Y(dp.rf._abc_6362_n7521) );
	NAND2X1 NAND2X1_5132 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7521), .Y(dp.rf._abc_6362_n7522) );
	NAND2X1 NAND2X1_5133 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<21>), .Y(dp.rf._abc_6362_n7523) );
	NAND2X1 NAND2X1_5134 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7523), .Y(dp.rf._abc_6362_n7524) );
	INVX1 INVX1_194 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<21>), .Y(dp.rf._abc_6362_n7525) );
	NOR2X1 NOR2X1_684 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7525), .Y(dp.rf._abc_6362_n7526) );
	NOR2X1 NOR2X1_685 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7524), .B(dp.rf._abc_6362_n7526), .Y(dp.rf._abc_6362_n7527) );
	NAND2X1 NAND2X1_5135 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<21>), .Y(dp.rf._abc_6362_n7528) );
	NAND2X1 NAND2X1_5136 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7528), .Y(dp.rf._abc_6362_n7529) );
	INVX1 INVX1_195 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<21>), .Y(dp.rf._abc_6362_n7530) );
	NOR2X1 NOR2X1_686 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7530), .Y(dp.rf._abc_6362_n7531) );
	NOR2X1 NOR2X1_687 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7529), .B(dp.rf._abc_6362_n7531), .Y(dp.rf._abc_6362_n7532) );
	OR2X2 OR2X2_65 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7527), .B(dp.rf._abc_6362_n7532), .Y(dp.rf._abc_6362_n7533) );
	NAND2X1 NAND2X1_5137 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7533), .Y(dp.rf._abc_6362_n7534) );
	AND2X2 AND2X2_260 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7534), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7535) );
	NAND2X1 NAND2X1_5138 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7522), .B(dp.rf._abc_6362_n7535), .Y(dp.rf._abc_6362_n7536) );
	NAND2X1 NAND2X1_5139 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<21>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7537) );
	NAND2X1 NAND2X1_5140 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<21>), .Y(dp.rf._abc_6362_n7538) );
	AND2X2 AND2X2_261 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7538), .B(instr[22]), .Y(dp.rf._abc_6362_n7539) );
	NAND2X1 NAND2X1_5141 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7537), .B(dp.rf._abc_6362_n7539), .Y(dp.rf._abc_6362_n7540) );
	NAND2X1 NAND2X1_5142 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<21>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7541) );
	NAND2X1 NAND2X1_5143 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<21>), .Y(dp.rf._abc_6362_n7542) );
	AND2X2 AND2X2_262 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7542), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7543) );
	NAND2X1 NAND2X1_5144 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7541), .B(dp.rf._abc_6362_n7543), .Y(dp.rf._abc_6362_n7544) );
	NAND2X1 NAND2X1_5145 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7540), .B(dp.rf._abc_6362_n7544), .Y(dp.rf._abc_6362_n7545) );
	AND2X2 AND2X2_263 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7545), .B(instr[23]), .Y(dp.rf._abc_6362_n7546) );
	NAND2X1 NAND2X1_5146 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<21>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7547) );
	NAND2X1 NAND2X1_5147 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<21>), .Y(dp.rf._abc_6362_n7548) );
	AND2X2 AND2X2_264 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7548), .B(instr[22]), .Y(dp.rf._abc_6362_n7549) );
	NAND2X1 NAND2X1_5148 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7547), .B(dp.rf._abc_6362_n7549), .Y(dp.rf._abc_6362_n7550) );
	NAND2X1 NAND2X1_5149 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<21>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7551) );
	NAND2X1 NAND2X1_5150 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<21>), .Y(dp.rf._abc_6362_n7552) );
	AND2X2 AND2X2_265 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7552), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7553) );
	NAND2X1 NAND2X1_5151 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7551), .B(dp.rf._abc_6362_n7553), .Y(dp.rf._abc_6362_n7554) );
	NAND2X1 NAND2X1_5152 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7550), .B(dp.rf._abc_6362_n7554), .Y(dp.rf._abc_6362_n7555) );
	NAND2X1 NAND2X1_5153 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7555), .Y(dp.rf._abc_6362_n7556) );
	NAND2X1 NAND2X1_5154 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7556), .Y(dp.rf._abc_6362_n7557) );
	NOR2X1 NOR2X1_688 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7546), .B(dp.rf._abc_6362_n7557), .Y(dp.rf._abc_6362_n7558) );
	NOR2X1 NOR2X1_689 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7558), .Y(dp.rf._abc_6362_n7559) );
	NAND2X1 NAND2X1_5155 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7536), .B(dp.rf._abc_6362_n7559), .Y(dp.rf._abc_6362_n7560) );
	NAND2X1 NAND2X1_5156 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n7560), .Y(dp.rf._abc_6362_n7561) );
	NOR2X1 NOR2X1_690 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7510), .B(dp.rf._abc_6362_n7561), .Y(dp.srca_21_) );
	NAND2X1 NAND2X1_5157 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<22>), .Y(dp.rf._abc_6362_n7563) );
	NAND2X1 NAND2X1_5158 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7563), .Y(dp.rf._abc_6362_n7564) );
	INVX1 INVX1_196 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<22>), .Y(dp.rf._abc_6362_n7565) );
	NOR2X1 NOR2X1_691 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7565), .Y(dp.rf._abc_6362_n7566) );
	NOR2X1 NOR2X1_692 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7564), .B(dp.rf._abc_6362_n7566), .Y(dp.rf._abc_6362_n7567) );
	NAND2X1 NAND2X1_5159 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<22>), .Y(dp.rf._abc_6362_n7568) );
	NAND2X1 NAND2X1_5160 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7568), .Y(dp.rf._abc_6362_n7569) );
	INVX1 INVX1_197 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<22>), .Y(dp.rf._abc_6362_n7570) );
	NOR2X1 NOR2X1_693 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7570), .Y(dp.rf._abc_6362_n7571) );
	NOR2X1 NOR2X1_694 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7569), .B(dp.rf._abc_6362_n7571), .Y(dp.rf._abc_6362_n7572) );
	NOR2X1 NOR2X1_695 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7567), .B(dp.rf._abc_6362_n7572), .Y(dp.rf._abc_6362_n7573) );
	NAND2X1 NAND2X1_5161 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7573), .Y(dp.rf._abc_6362_n7574) );
	NAND2X1 NAND2X1_5162 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<22>), .Y(dp.rf._abc_6362_n7575) );
	NAND2X1 NAND2X1_5163 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7575), .Y(dp.rf._abc_6362_n7576) );
	INVX1 INVX1_198 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<22>), .Y(dp.rf._abc_6362_n7577) );
	NOR2X1 NOR2X1_696 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7577), .Y(dp.rf._abc_6362_n7578) );
	NOR2X1 NOR2X1_697 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7576), .B(dp.rf._abc_6362_n7578), .Y(dp.rf._abc_6362_n7579) );
	NAND2X1 NAND2X1_5164 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<22>), .Y(dp.rf._abc_6362_n7580) );
	NAND2X1 NAND2X1_5165 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7580), .Y(dp.rf._abc_6362_n7581) );
	INVX1 INVX1_199 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<22>), .Y(dp.rf._abc_6362_n7582) );
	NOR2X1 NOR2X1_698 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7582), .Y(dp.rf._abc_6362_n7583) );
	NOR2X1 NOR2X1_699 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7581), .B(dp.rf._abc_6362_n7583), .Y(dp.rf._abc_6362_n7584) );
	NOR2X1 NOR2X1_700 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7579), .B(dp.rf._abc_6362_n7584), .Y(dp.rf._abc_6362_n7585) );
	NAND2X1 NAND2X1_5166 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7585), .Y(dp.rf._abc_6362_n7586) );
	NAND2X1 NAND2X1_5167 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7574), .B(dp.rf._abc_6362_n7586), .Y(dp.rf._abc_6362_n7587) );
	NAND2X1 NAND2X1_5168 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7587), .Y(dp.rf._abc_6362_n7588) );
	NAND2X1 NAND2X1_5169 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7588), .Y(dp.rf._abc_6362_n7589) );
	NAND2X1 NAND2X1_5170 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<22>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7590) );
	INVX1 INVX1_200 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<22>), .Y(dp.rf._abc_6362_n7591) );
	NOR2X1 NOR2X1_701 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7591), .Y(dp.rf._abc_6362_n7592) );
	NOR2X1 NOR2X1_702 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7592), .Y(dp.rf._abc_6362_n7593) );
	NAND2X1 NAND2X1_5171 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7590), .B(dp.rf._abc_6362_n7593), .Y(dp.rf._abc_6362_n7594) );
	NAND2X1 NAND2X1_5172 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<22>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7595) );
	INVX1 INVX1_201 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<22>), .Y(dp.rf._abc_6362_n7596) );
	NOR2X1 NOR2X1_703 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7596), .Y(dp.rf._abc_6362_n7597) );
	NOR2X1 NOR2X1_704 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7597), .Y(dp.rf._abc_6362_n7598) );
	NAND2X1 NAND2X1_5173 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7595), .B(dp.rf._abc_6362_n7598), .Y(dp.rf._abc_6362_n7599) );
	NAND2X1 NAND2X1_5174 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7594), .B(dp.rf._abc_6362_n7599), .Y(dp.rf._abc_6362_n7600) );
	NOR2X1 NOR2X1_705 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7600), .Y(dp.rf._abc_6362_n7601) );
	NAND2X1 NAND2X1_5175 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<22>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7602) );
	INVX1 INVX1_202 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<22>), .Y(dp.rf._abc_6362_n7603) );
	NOR2X1 NOR2X1_706 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7603), .Y(dp.rf._abc_6362_n7604) );
	NOR2X1 NOR2X1_707 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7604), .Y(dp.rf._abc_6362_n7605) );
	NAND2X1 NAND2X1_5176 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7602), .B(dp.rf._abc_6362_n7605), .Y(dp.rf._abc_6362_n7606) );
	NAND2X1 NAND2X1_5177 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<22>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7607) );
	INVX1 INVX1_203 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<22>), .Y(dp.rf._abc_6362_n7608) );
	NOR2X1 NOR2X1_708 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7608), .Y(dp.rf._abc_6362_n7609) );
	NOR2X1 NOR2X1_709 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7609), .Y(dp.rf._abc_6362_n7610) );
	NAND2X1 NAND2X1_5178 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7607), .B(dp.rf._abc_6362_n7610), .Y(dp.rf._abc_6362_n7611) );
	NAND2X1 NAND2X1_5179 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7606), .B(dp.rf._abc_6362_n7611), .Y(dp.rf._abc_6362_n7612) );
	NOR2X1 NOR2X1_710 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7612), .Y(dp.rf._abc_6362_n7613) );
	NOR2X1 NOR2X1_711 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7601), .B(dp.rf._abc_6362_n7613), .Y(dp.rf._abc_6362_n7614) );
	NOR2X1 NOR2X1_712 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7614), .Y(dp.rf._abc_6362_n7615) );
	NOR2X1 NOR2X1_713 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7589), .B(dp.rf._abc_6362_n7615), .Y(dp.rf._abc_6362_n7616) );
	NAND2X1 NAND2X1_5180 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<22>), .Y(dp.rf._abc_6362_n7617) );
	NAND2X1 NAND2X1_5181 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7617), .Y(dp.rf._abc_6362_n7618) );
	INVX1 INVX1_204 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<22>), .Y(dp.rf._abc_6362_n7619) );
	NOR2X1 NOR2X1_714 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7619), .Y(dp.rf._abc_6362_n7620) );
	NOR2X1 NOR2X1_715 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7618), .B(dp.rf._abc_6362_n7620), .Y(dp.rf._abc_6362_n7621) );
	NAND2X1 NAND2X1_5182 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<22>), .Y(dp.rf._abc_6362_n7622) );
	NAND2X1 NAND2X1_5183 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7622), .Y(dp.rf._abc_6362_n7623) );
	INVX1 INVX1_205 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<22>), .Y(dp.rf._abc_6362_n7624) );
	NOR2X1 NOR2X1_716 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7624), .Y(dp.rf._abc_6362_n7625) );
	NOR2X1 NOR2X1_717 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7623), .B(dp.rf._abc_6362_n7625), .Y(dp.rf._abc_6362_n7626) );
	OR2X2 OR2X2_66 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7621), .B(dp.rf._abc_6362_n7626), .Y(dp.rf._abc_6362_n7627) );
	NAND2X1 NAND2X1_5184 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7627), .Y(dp.rf._abc_6362_n7628) );
	NAND2X1 NAND2X1_5185 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<22>), .Y(dp.rf._abc_6362_n7629) );
	NAND2X1 NAND2X1_5186 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7629), .Y(dp.rf._abc_6362_n7630) );
	INVX1 INVX1_206 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<22>), .Y(dp.rf._abc_6362_n7631) );
	NOR2X1 NOR2X1_718 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7631), .Y(dp.rf._abc_6362_n7632) );
	NOR2X1 NOR2X1_719 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7630), .B(dp.rf._abc_6362_n7632), .Y(dp.rf._abc_6362_n7633) );
	NAND2X1 NAND2X1_5187 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<22>), .Y(dp.rf._abc_6362_n7634) );
	NAND2X1 NAND2X1_5188 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7634), .Y(dp.rf._abc_6362_n7635) );
	INVX1 INVX1_207 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<22>), .Y(dp.rf._abc_6362_n7636) );
	NOR2X1 NOR2X1_720 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7636), .Y(dp.rf._abc_6362_n7637) );
	NOR2X1 NOR2X1_721 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7635), .B(dp.rf._abc_6362_n7637), .Y(dp.rf._abc_6362_n7638) );
	OR2X2 OR2X2_67 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7633), .B(dp.rf._abc_6362_n7638), .Y(dp.rf._abc_6362_n7639) );
	NAND2X1 NAND2X1_5189 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7639), .Y(dp.rf._abc_6362_n7640) );
	AND2X2 AND2X2_266 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7640), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7641) );
	NAND2X1 NAND2X1_5190 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7628), .B(dp.rf._abc_6362_n7641), .Y(dp.rf._abc_6362_n7642) );
	NAND2X1 NAND2X1_5191 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<22>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7643) );
	NAND2X1 NAND2X1_5192 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<22>), .Y(dp.rf._abc_6362_n7644) );
	AND2X2 AND2X2_267 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7644), .B(instr[22]), .Y(dp.rf._abc_6362_n7645) );
	NAND2X1 NAND2X1_5193 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7643), .B(dp.rf._abc_6362_n7645), .Y(dp.rf._abc_6362_n7646) );
	NAND2X1 NAND2X1_5194 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<22>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7647) );
	NAND2X1 NAND2X1_5195 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<22>), .Y(dp.rf._abc_6362_n7648) );
	AND2X2 AND2X2_268 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7648), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7649) );
	NAND2X1 NAND2X1_5196 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7647), .B(dp.rf._abc_6362_n7649), .Y(dp.rf._abc_6362_n7650) );
	NAND2X1 NAND2X1_5197 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7646), .B(dp.rf._abc_6362_n7650), .Y(dp.rf._abc_6362_n7651) );
	AND2X2 AND2X2_269 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7651), .B(instr[23]), .Y(dp.rf._abc_6362_n7652) );
	NAND2X1 NAND2X1_5198 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<22>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7653) );
	NAND2X1 NAND2X1_5199 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<22>), .Y(dp.rf._abc_6362_n7654) );
	AND2X2 AND2X2_270 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7654), .B(instr[22]), .Y(dp.rf._abc_6362_n7655) );
	NAND2X1 NAND2X1_5200 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7653), .B(dp.rf._abc_6362_n7655), .Y(dp.rf._abc_6362_n7656) );
	NAND2X1 NAND2X1_5201 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<22>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7657) );
	NAND2X1 NAND2X1_5202 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<22>), .Y(dp.rf._abc_6362_n7658) );
	AND2X2 AND2X2_271 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7658), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7659) );
	NAND2X1 NAND2X1_5203 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7657), .B(dp.rf._abc_6362_n7659), .Y(dp.rf._abc_6362_n7660) );
	NAND2X1 NAND2X1_5204 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7656), .B(dp.rf._abc_6362_n7660), .Y(dp.rf._abc_6362_n7661) );
	NAND2X1 NAND2X1_5205 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7661), .Y(dp.rf._abc_6362_n7662) );
	NAND2X1 NAND2X1_5206 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7662), .Y(dp.rf._abc_6362_n7663) );
	NOR2X1 NOR2X1_722 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7652), .B(dp.rf._abc_6362_n7663), .Y(dp.rf._abc_6362_n7664) );
	NOR2X1 NOR2X1_723 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7664), .Y(dp.rf._abc_6362_n7665) );
	NAND2X1 NAND2X1_5207 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7642), .B(dp.rf._abc_6362_n7665), .Y(dp.rf._abc_6362_n7666) );
	NAND2X1 NAND2X1_5208 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n7666), .Y(dp.rf._abc_6362_n7667) );
	NOR2X1 NOR2X1_724 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7616), .B(dp.rf._abc_6362_n7667), .Y(dp.srca_22_) );
	NAND2X1 NAND2X1_5209 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<23>), .Y(dp.rf._abc_6362_n7669) );
	NAND2X1 NAND2X1_5210 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7669), .Y(dp.rf._abc_6362_n7670) );
	INVX1 INVX1_208 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<23>), .Y(dp.rf._abc_6362_n7671) );
	NOR2X1 NOR2X1_725 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7671), .Y(dp.rf._abc_6362_n7672) );
	NOR2X1 NOR2X1_726 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7670), .B(dp.rf._abc_6362_n7672), .Y(dp.rf._abc_6362_n7673) );
	NAND2X1 NAND2X1_5211 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<23>), .Y(dp.rf._abc_6362_n7674) );
	NAND2X1 NAND2X1_5212 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7674), .Y(dp.rf._abc_6362_n7675) );
	INVX1 INVX1_209 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<23>), .Y(dp.rf._abc_6362_n7676) );
	NOR2X1 NOR2X1_727 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7676), .Y(dp.rf._abc_6362_n7677) );
	NOR2X1 NOR2X1_728 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7675), .B(dp.rf._abc_6362_n7677), .Y(dp.rf._abc_6362_n7678) );
	NOR2X1 NOR2X1_729 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7673), .B(dp.rf._abc_6362_n7678), .Y(dp.rf._abc_6362_n7679) );
	NAND2X1 NAND2X1_5213 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7679), .Y(dp.rf._abc_6362_n7680) );
	NAND2X1 NAND2X1_5214 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<23>), .Y(dp.rf._abc_6362_n7681) );
	NAND2X1 NAND2X1_5215 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7681), .Y(dp.rf._abc_6362_n7682) );
	INVX1 INVX1_210 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<23>), .Y(dp.rf._abc_6362_n7683) );
	NOR2X1 NOR2X1_730 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7683), .Y(dp.rf._abc_6362_n7684) );
	NOR2X1 NOR2X1_731 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7682), .B(dp.rf._abc_6362_n7684), .Y(dp.rf._abc_6362_n7685) );
	NAND2X1 NAND2X1_5216 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<23>), .Y(dp.rf._abc_6362_n7686) );
	NAND2X1 NAND2X1_5217 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7686), .Y(dp.rf._abc_6362_n7687) );
	INVX1 INVX1_211 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<23>), .Y(dp.rf._abc_6362_n7688) );
	NOR2X1 NOR2X1_732 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7688), .Y(dp.rf._abc_6362_n7689) );
	NOR2X1 NOR2X1_733 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7687), .B(dp.rf._abc_6362_n7689), .Y(dp.rf._abc_6362_n7690) );
	NOR2X1 NOR2X1_734 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7685), .B(dp.rf._abc_6362_n7690), .Y(dp.rf._abc_6362_n7691) );
	NAND2X1 NAND2X1_5218 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7691), .Y(dp.rf._abc_6362_n7692) );
	NAND2X1 NAND2X1_5219 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7680), .B(dp.rf._abc_6362_n7692), .Y(dp.rf._abc_6362_n7693) );
	NAND2X1 NAND2X1_5220 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7693), .Y(dp.rf._abc_6362_n7694) );
	NAND2X1 NAND2X1_5221 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7694), .Y(dp.rf._abc_6362_n7695) );
	NAND2X1 NAND2X1_5222 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7696) );
	INVX1 INVX1_212 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<23>), .Y(dp.rf._abc_6362_n7697) );
	NOR2X1 NOR2X1_735 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7697), .Y(dp.rf._abc_6362_n7698) );
	NOR2X1 NOR2X1_736 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7698), .Y(dp.rf._abc_6362_n7699) );
	NAND2X1 NAND2X1_5223 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7696), .B(dp.rf._abc_6362_n7699), .Y(dp.rf._abc_6362_n7700) );
	NAND2X1 NAND2X1_5224 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7701) );
	INVX1 INVX1_213 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<23>), .Y(dp.rf._abc_6362_n7702) );
	NOR2X1 NOR2X1_737 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7702), .Y(dp.rf._abc_6362_n7703) );
	NOR2X1 NOR2X1_738 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7703), .Y(dp.rf._abc_6362_n7704) );
	NAND2X1 NAND2X1_5225 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7701), .B(dp.rf._abc_6362_n7704), .Y(dp.rf._abc_6362_n7705) );
	NAND2X1 NAND2X1_5226 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7700), .B(dp.rf._abc_6362_n7705), .Y(dp.rf._abc_6362_n7706) );
	NOR2X1 NOR2X1_739 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7706), .Y(dp.rf._abc_6362_n7707) );
	NAND2X1 NAND2X1_5227 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7708) );
	INVX1 INVX1_214 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<23>), .Y(dp.rf._abc_6362_n7709) );
	NOR2X1 NOR2X1_740 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7709), .Y(dp.rf._abc_6362_n7710) );
	NOR2X1 NOR2X1_741 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7710), .Y(dp.rf._abc_6362_n7711) );
	NAND2X1 NAND2X1_5228 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7708), .B(dp.rf._abc_6362_n7711), .Y(dp.rf._abc_6362_n7712) );
	NAND2X1 NAND2X1_5229 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7713) );
	INVX1 INVX1_215 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<23>), .Y(dp.rf._abc_6362_n7714) );
	NOR2X1 NOR2X1_742 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7714), .Y(dp.rf._abc_6362_n7715) );
	NOR2X1 NOR2X1_743 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7715), .Y(dp.rf._abc_6362_n7716) );
	NAND2X1 NAND2X1_5230 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7713), .B(dp.rf._abc_6362_n7716), .Y(dp.rf._abc_6362_n7717) );
	NAND2X1 NAND2X1_5231 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7712), .B(dp.rf._abc_6362_n7717), .Y(dp.rf._abc_6362_n7718) );
	NOR2X1 NOR2X1_744 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7718), .Y(dp.rf._abc_6362_n7719) );
	NOR2X1 NOR2X1_745 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7707), .B(dp.rf._abc_6362_n7719), .Y(dp.rf._abc_6362_n7720) );
	NOR2X1 NOR2X1_746 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7720), .Y(dp.rf._abc_6362_n7721) );
	NOR2X1 NOR2X1_747 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7695), .B(dp.rf._abc_6362_n7721), .Y(dp.rf._abc_6362_n7722) );
	NAND2X1 NAND2X1_5232 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<23>), .Y(dp.rf._abc_6362_n7723) );
	NAND2X1 NAND2X1_5233 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7724) );
	NAND2X1 NAND2X1_5234 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7723), .B(dp.rf._abc_6362_n7724), .Y(dp.rf._abc_6362_n7725) );
	NAND2X1 NAND2X1_5235 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7725), .Y(dp.rf._abc_6362_n7726) );
	NAND2X1 NAND2X1_5236 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<23>), .Y(dp.rf._abc_6362_n7727) );
	NAND2X1 NAND2X1_5237 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7728) );
	NAND2X1 NAND2X1_5238 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7727), .B(dp.rf._abc_6362_n7728), .Y(dp.rf._abc_6362_n7729) );
	NAND2X1 NAND2X1_5239 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7729), .Y(dp.rf._abc_6362_n7730) );
	AND2X2 AND2X2_272 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7726), .B(dp.rf._abc_6362_n7730), .Y(dp.rf._abc_6362_n7731) );
	NAND2X1 NAND2X1_5240 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7731), .Y(dp.rf._abc_6362_n7732) );
	NAND2X1 NAND2X1_5241 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<23>), .Y(dp.rf._abc_6362_n7733) );
	NAND2X1 NAND2X1_5242 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7734) );
	NAND2X1 NAND2X1_5243 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7733), .B(dp.rf._abc_6362_n7734), .Y(dp.rf._abc_6362_n7735) );
	NAND2X1 NAND2X1_5244 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7735), .Y(dp.rf._abc_6362_n7736) );
	NAND2X1 NAND2X1_5245 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<23>), .Y(dp.rf._abc_6362_n7737) );
	NAND2X1 NAND2X1_5246 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7738) );
	NAND2X1 NAND2X1_5247 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7737), .B(dp.rf._abc_6362_n7738), .Y(dp.rf._abc_6362_n7739) );
	NAND2X1 NAND2X1_5248 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7739), .Y(dp.rf._abc_6362_n7740) );
	AND2X2 AND2X2_273 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7736), .B(dp.rf._abc_6362_n7740), .Y(dp.rf._abc_6362_n7741) );
	NAND2X1 NAND2X1_5249 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7741), .Y(dp.rf._abc_6362_n7742) );
	AND2X2 AND2X2_274 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7742), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7743) );
	NAND2X1 NAND2X1_5250 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7732), .B(dp.rf._abc_6362_n7743), .Y(dp.rf._abc_6362_n7744) );
	NAND2X1 NAND2X1_5251 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7745) );
	NAND2X1 NAND2X1_5252 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<23>), .Y(dp.rf._abc_6362_n7746) );
	AND2X2 AND2X2_275 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7746), .B(instr[22]), .Y(dp.rf._abc_6362_n7747) );
	NAND2X1 NAND2X1_5253 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7745), .B(dp.rf._abc_6362_n7747), .Y(dp.rf._abc_6362_n7748) );
	NAND2X1 NAND2X1_5254 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7749) );
	NAND2X1 NAND2X1_5255 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<23>), .Y(dp.rf._abc_6362_n7750) );
	AND2X2 AND2X2_276 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7750), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7751) );
	NAND2X1 NAND2X1_5256 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7749), .B(dp.rf._abc_6362_n7751), .Y(dp.rf._abc_6362_n7752) );
	NAND2X1 NAND2X1_5257 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7748), .B(dp.rf._abc_6362_n7752), .Y(dp.rf._abc_6362_n7753) );
	AND2X2 AND2X2_277 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7753), .B(instr[23]), .Y(dp.rf._abc_6362_n7754) );
	NAND2X1 NAND2X1_5258 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7755) );
	NAND2X1 NAND2X1_5259 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<23>), .Y(dp.rf._abc_6362_n7756) );
	AND2X2 AND2X2_278 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7756), .B(instr[22]), .Y(dp.rf._abc_6362_n7757) );
	NAND2X1 NAND2X1_5260 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7755), .B(dp.rf._abc_6362_n7757), .Y(dp.rf._abc_6362_n7758) );
	NAND2X1 NAND2X1_5261 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<23>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7759) );
	NAND2X1 NAND2X1_5262 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<23>), .Y(dp.rf._abc_6362_n7760) );
	AND2X2 AND2X2_279 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7760), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7761) );
	NAND2X1 NAND2X1_5263 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7759), .B(dp.rf._abc_6362_n7761), .Y(dp.rf._abc_6362_n7762) );
	NAND2X1 NAND2X1_5264 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7758), .B(dp.rf._abc_6362_n7762), .Y(dp.rf._abc_6362_n7763) );
	NAND2X1 NAND2X1_5265 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7763), .Y(dp.rf._abc_6362_n7764) );
	NAND2X1 NAND2X1_5266 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7764), .Y(dp.rf._abc_6362_n7765) );
	NOR2X1 NOR2X1_748 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7754), .B(dp.rf._abc_6362_n7765), .Y(dp.rf._abc_6362_n7766) );
	NOR2X1 NOR2X1_749 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7766), .Y(dp.rf._abc_6362_n7767) );
	NAND2X1 NAND2X1_5267 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7744), .B(dp.rf._abc_6362_n7767), .Y(dp.rf._abc_6362_n7768) );
	NAND2X1 NAND2X1_5268 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n7768), .Y(dp.rf._abc_6362_n7769) );
	NOR2X1 NOR2X1_750 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7722), .B(dp.rf._abc_6362_n7769), .Y(dp.srca_23_) );
	NAND2X1 NAND2X1_5269 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7771) );
	INVX1 INVX1_216 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<24>), .Y(dp.rf._abc_6362_n7772) );
	NOR2X1 NOR2X1_751 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7772), .Y(dp.rf._abc_6362_n7773) );
	NOR2X1 NOR2X1_752 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7773), .Y(dp.rf._abc_6362_n7774) );
	NAND2X1 NAND2X1_5270 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7771), .B(dp.rf._abc_6362_n7774), .Y(dp.rf._abc_6362_n7775) );
	NAND2X1 NAND2X1_5271 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7776) );
	INVX1 INVX1_217 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<24>), .Y(dp.rf._abc_6362_n7777) );
	NOR2X1 NOR2X1_753 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7777), .Y(dp.rf._abc_6362_n7778) );
	NOR2X1 NOR2X1_754 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7778), .Y(dp.rf._abc_6362_n7779) );
	NAND2X1 NAND2X1_5272 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7776), .B(dp.rf._abc_6362_n7779), .Y(dp.rf._abc_6362_n7780) );
	NAND2X1 NAND2X1_5273 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7775), .B(dp.rf._abc_6362_n7780), .Y(dp.rf._abc_6362_n7781) );
	NAND2X1 NAND2X1_5274 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7781), .Y(dp.rf._abc_6362_n7782) );
	NAND2X1 NAND2X1_5275 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7783) );
	INVX1 INVX1_218 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<24>), .Y(dp.rf._abc_6362_n7784) );
	NOR2X1 NOR2X1_755 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7784), .Y(dp.rf._abc_6362_n7785) );
	NOR2X1 NOR2X1_756 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7785), .Y(dp.rf._abc_6362_n7786) );
	NAND2X1 NAND2X1_5276 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7783), .B(dp.rf._abc_6362_n7786), .Y(dp.rf._abc_6362_n7787) );
	NAND2X1 NAND2X1_5277 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7788) );
	INVX1 INVX1_219 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<24>), .Y(dp.rf._abc_6362_n7789) );
	NOR2X1 NOR2X1_757 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7789), .Y(dp.rf._abc_6362_n7790) );
	NOR2X1 NOR2X1_758 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7790), .Y(dp.rf._abc_6362_n7791) );
	NAND2X1 NAND2X1_5278 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7788), .B(dp.rf._abc_6362_n7791), .Y(dp.rf._abc_6362_n7792) );
	NAND2X1 NAND2X1_5279 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7787), .B(dp.rf._abc_6362_n7792), .Y(dp.rf._abc_6362_n7793) );
	NAND2X1 NAND2X1_5280 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7793), .Y(dp.rf._abc_6362_n7794) );
	NAND2X1 NAND2X1_5281 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7782), .B(dp.rf._abc_6362_n7794), .Y(dp.rf._abc_6362_n7795) );
	NOR2X1 NOR2X1_759 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7795), .Y(dp.rf._abc_6362_n7796) );
	NAND2X1 NAND2X1_5282 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<24>), .Y(dp.rf._abc_6362_n7797) );
	NAND2X1 NAND2X1_5283 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7797), .Y(dp.rf._abc_6362_n7798) );
	INVX1 INVX1_220 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<24>), .Y(dp.rf._abc_6362_n7799) );
	NOR2X1 NOR2X1_760 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7799), .Y(dp.rf._abc_6362_n7800) );
	NOR2X1 NOR2X1_761 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7798), .B(dp.rf._abc_6362_n7800), .Y(dp.rf._abc_6362_n7801) );
	NAND2X1 NAND2X1_5284 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<24>), .Y(dp.rf._abc_6362_n7802) );
	NAND2X1 NAND2X1_5285 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7802), .Y(dp.rf._abc_6362_n7803) );
	INVX1 INVX1_221 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<24>), .Y(dp.rf._abc_6362_n7804) );
	NOR2X1 NOR2X1_762 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7804), .Y(dp.rf._abc_6362_n7805) );
	NOR2X1 NOR2X1_763 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7803), .B(dp.rf._abc_6362_n7805), .Y(dp.rf._abc_6362_n7806) );
	OR2X2 OR2X2_68 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7801), .B(dp.rf._abc_6362_n7806), .Y(dp.rf._abc_6362_n7807) );
	NAND2X1 NAND2X1_5286 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7807), .Y(dp.rf._abc_6362_n7808) );
	NAND2X1 NAND2X1_5287 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<24>), .Y(dp.rf._abc_6362_n7809) );
	NAND2X1 NAND2X1_5288 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7809), .Y(dp.rf._abc_6362_n7810) );
	INVX1 INVX1_222 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<24>), .Y(dp.rf._abc_6362_n7811) );
	NOR2X1 NOR2X1_764 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7811), .Y(dp.rf._abc_6362_n7812) );
	NOR2X1 NOR2X1_765 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7810), .B(dp.rf._abc_6362_n7812), .Y(dp.rf._abc_6362_n7813) );
	NAND2X1 NAND2X1_5289 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<24>), .Y(dp.rf._abc_6362_n7814) );
	NAND2X1 NAND2X1_5290 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7814), .Y(dp.rf._abc_6362_n7815) );
	INVX1 INVX1_223 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<24>), .Y(dp.rf._abc_6362_n7816) );
	NOR2X1 NOR2X1_766 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7816), .Y(dp.rf._abc_6362_n7817) );
	NOR2X1 NOR2X1_767 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7815), .B(dp.rf._abc_6362_n7817), .Y(dp.rf._abc_6362_n7818) );
	OR2X2 OR2X2_69 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7813), .B(dp.rf._abc_6362_n7818), .Y(dp.rf._abc_6362_n7819) );
	NAND2X1 NAND2X1_5291 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7819), .Y(dp.rf._abc_6362_n7820) );
	AND2X2 AND2X2_280 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7820), .B(instr[24]), .Y(dp.rf._abc_6362_n7821) );
	NAND2X1 NAND2X1_5292 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7808), .B(dp.rf._abc_6362_n7821), .Y(dp.rf._abc_6362_n7822) );
	NAND2X1 NAND2X1_5293 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7822), .Y(dp.rf._abc_6362_n7823) );
	NOR2X1 NOR2X1_768 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7796), .B(dp.rf._abc_6362_n7823), .Y(dp.rf._abc_6362_n7824) );
	NAND2X1 NAND2X1_5294 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<24>), .Y(dp.rf._abc_6362_n7825) );
	NAND2X1 NAND2X1_5295 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7826) );
	NAND2X1 NAND2X1_5296 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7825), .B(dp.rf._abc_6362_n7826), .Y(dp.rf._abc_6362_n7827) );
	NAND2X1 NAND2X1_5297 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7827), .Y(dp.rf._abc_6362_n7828) );
	NAND2X1 NAND2X1_5298 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<24>), .Y(dp.rf._abc_6362_n7829) );
	NAND2X1 NAND2X1_5299 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7830) );
	NAND2X1 NAND2X1_5300 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7829), .B(dp.rf._abc_6362_n7830), .Y(dp.rf._abc_6362_n7831) );
	NAND2X1 NAND2X1_5301 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7831), .Y(dp.rf._abc_6362_n7832) );
	NAND2X1 NAND2X1_5302 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7828), .B(dp.rf._abc_6362_n7832), .Y(dp.rf._abc_6362_n7833) );
	NAND2X1 NAND2X1_5303 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7833), .Y(dp.rf._abc_6362_n7834) );
	NAND2X1 NAND2X1_5304 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<24>), .Y(dp.rf._abc_6362_n7835) );
	NAND2X1 NAND2X1_5305 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7836) );
	NAND2X1 NAND2X1_5306 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7835), .B(dp.rf._abc_6362_n7836), .Y(dp.rf._abc_6362_n7837) );
	NAND2X1 NAND2X1_5307 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7837), .Y(dp.rf._abc_6362_n7838) );
	NAND2X1 NAND2X1_5308 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<24>), .Y(dp.rf._abc_6362_n7839) );
	NAND2X1 NAND2X1_5309 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7840) );
	NAND2X1 NAND2X1_5310 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7839), .B(dp.rf._abc_6362_n7840), .Y(dp.rf._abc_6362_n7841) );
	NAND2X1 NAND2X1_5311 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7841), .Y(dp.rf._abc_6362_n7842) );
	NAND2X1 NAND2X1_5312 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7838), .B(dp.rf._abc_6362_n7842), .Y(dp.rf._abc_6362_n7843) );
	NAND2X1 NAND2X1_5313 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7843), .Y(dp.rf._abc_6362_n7844) );
	NAND2X1 NAND2X1_5314 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7834), .B(dp.rf._abc_6362_n7844), .Y(dp.rf._abc_6362_n7845) );
	NAND2X1 NAND2X1_5315 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7845), .Y(dp.rf._abc_6362_n7846) );
	NAND2X1 NAND2X1_5316 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7847) );
	NAND2X1 NAND2X1_5317 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<24>), .Y(dp.rf._abc_6362_n7848) );
	AND2X2 AND2X2_281 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7848), .B(instr[22]), .Y(dp.rf._abc_6362_n7849) );
	NAND2X1 NAND2X1_5318 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7847), .B(dp.rf._abc_6362_n7849), .Y(dp.rf._abc_6362_n7850) );
	NAND2X1 NAND2X1_5319 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7851) );
	NAND2X1 NAND2X1_5320 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<24>), .Y(dp.rf._abc_6362_n7852) );
	AND2X2 AND2X2_282 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7852), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7853) );
	NAND2X1 NAND2X1_5321 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7851), .B(dp.rf._abc_6362_n7853), .Y(dp.rf._abc_6362_n7854) );
	NAND2X1 NAND2X1_5322 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7850), .B(dp.rf._abc_6362_n7854), .Y(dp.rf._abc_6362_n7855) );
	AND2X2 AND2X2_283 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7855), .B(instr[23]), .Y(dp.rf._abc_6362_n7856) );
	NAND2X1 NAND2X1_5323 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7857) );
	NAND2X1 NAND2X1_5324 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<24>), .Y(dp.rf._abc_6362_n7858) );
	AND2X2 AND2X2_284 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7858), .B(instr[22]), .Y(dp.rf._abc_6362_n7859) );
	NAND2X1 NAND2X1_5325 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7857), .B(dp.rf._abc_6362_n7859), .Y(dp.rf._abc_6362_n7860) );
	NAND2X1 NAND2X1_5326 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<24>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7861) );
	NAND2X1 NAND2X1_5327 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<24>), .Y(dp.rf._abc_6362_n7862) );
	AND2X2 AND2X2_285 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7862), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7863) );
	NAND2X1 NAND2X1_5328 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7861), .B(dp.rf._abc_6362_n7863), .Y(dp.rf._abc_6362_n7864) );
	NAND2X1 NAND2X1_5329 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7860), .B(dp.rf._abc_6362_n7864), .Y(dp.rf._abc_6362_n7865) );
	NAND2X1 NAND2X1_5330 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7865), .Y(dp.rf._abc_6362_n7866) );
	NAND2X1 NAND2X1_5331 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n7866), .Y(dp.rf._abc_6362_n7867) );
	NOR2X1 NOR2X1_769 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7856), .B(dp.rf._abc_6362_n7867), .Y(dp.rf._abc_6362_n7868) );
	NOR2X1 NOR2X1_770 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7868), .Y(dp.rf._abc_6362_n7869) );
	NAND2X1 NAND2X1_5332 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7846), .B(dp.rf._abc_6362_n7869), .Y(dp.rf._abc_6362_n7870) );
	NAND2X1 NAND2X1_5333 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n7870), .Y(dp.rf._abc_6362_n7871) );
	NOR2X1 NOR2X1_771 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7824), .B(dp.rf._abc_6362_n7871), .Y(dp.srca_24_) );
	NAND2X1 NAND2X1_5334 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7873) );
	INVX1 INVX1_224 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_7_<25>), .Y(dp.rf._abc_6362_n7874) );
	NOR2X1 NOR2X1_772 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7874), .Y(dp.rf._abc_6362_n7875) );
	NOR2X1 NOR2X1_773 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7875), .Y(dp.rf._abc_6362_n7876) );
	NAND2X1 NAND2X1_5335 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7873), .B(dp.rf._abc_6362_n7876), .Y(dp.rf._abc_6362_n7877) );
	NAND2X1 NAND2X1_5336 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7878) );
	INVX1 INVX1_225 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_5_<25>), .Y(dp.rf._abc_6362_n7879) );
	NOR2X1 NOR2X1_774 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7879), .Y(dp.rf._abc_6362_n7880) );
	NOR2X1 NOR2X1_775 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7880), .Y(dp.rf._abc_6362_n7881) );
	NAND2X1 NAND2X1_5337 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7878), .B(dp.rf._abc_6362_n7881), .Y(dp.rf._abc_6362_n7882) );
	NAND2X1 NAND2X1_5338 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7877), .B(dp.rf._abc_6362_n7882), .Y(dp.rf._abc_6362_n7883) );
	NAND2X1 NAND2X1_5339 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7883), .Y(dp.rf._abc_6362_n7884) );
	NAND2X1 NAND2X1_5340 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7885) );
	INVX1 INVX1_226 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_3_<25>), .Y(dp.rf._abc_6362_n7886) );
	NOR2X1 NOR2X1_776 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7886), .Y(dp.rf._abc_6362_n7887) );
	NOR2X1 NOR2X1_777 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7887), .Y(dp.rf._abc_6362_n7888) );
	NAND2X1 NAND2X1_5341 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7885), .B(dp.rf._abc_6362_n7888), .Y(dp.rf._abc_6362_n7889) );
	NAND2X1 NAND2X1_5342 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7890) );
	INVX1 INVX1_227 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_1_<25>), .Y(dp.rf._abc_6362_n7891) );
	NOR2X1 NOR2X1_778 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf._abc_6362_n7891), .Y(dp.rf._abc_6362_n7892) );
	NOR2X1 NOR2X1_779 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7892), .Y(dp.rf._abc_6362_n7893) );
	NAND2X1 NAND2X1_5343 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7890), .B(dp.rf._abc_6362_n7893), .Y(dp.rf._abc_6362_n7894) );
	NAND2X1 NAND2X1_5344 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7889), .B(dp.rf._abc_6362_n7894), .Y(dp.rf._abc_6362_n7895) );
	NAND2X1 NAND2X1_5345 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7895), .Y(dp.rf._abc_6362_n7896) );
	NAND2X1 NAND2X1_5346 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7884), .B(dp.rf._abc_6362_n7896), .Y(dp.rf._abc_6362_n7897) );
	NOR2X1 NOR2X1_780 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7897), .Y(dp.rf._abc_6362_n7898) );
	NAND2X1 NAND2X1_5347 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<25>), .Y(dp.rf._abc_6362_n7899) );
	NAND2X1 NAND2X1_5348 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7899), .Y(dp.rf._abc_6362_n7900) );
	INVX1 INVX1_228 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<25>), .Y(dp.rf._abc_6362_n7901) );
	NOR2X1 NOR2X1_781 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7901), .Y(dp.rf._abc_6362_n7902) );
	NOR2X1 NOR2X1_782 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7900), .B(dp.rf._abc_6362_n7902), .Y(dp.rf._abc_6362_n7903) );
	NAND2X1 NAND2X1_5349 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<25>), .Y(dp.rf._abc_6362_n7904) );
	NAND2X1 NAND2X1_5350 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7904), .Y(dp.rf._abc_6362_n7905) );
	INVX1 INVX1_229 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<25>), .Y(dp.rf._abc_6362_n7906) );
	NOR2X1 NOR2X1_783 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7906), .Y(dp.rf._abc_6362_n7907) );
	NOR2X1 NOR2X1_784 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7905), .B(dp.rf._abc_6362_n7907), .Y(dp.rf._abc_6362_n7908) );
	OR2X2 OR2X2_70 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7903), .B(dp.rf._abc_6362_n7908), .Y(dp.rf._abc_6362_n7909) );
	NAND2X1 NAND2X1_5351 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7909), .Y(dp.rf._abc_6362_n7910) );
	NAND2X1 NAND2X1_5352 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<25>), .Y(dp.rf._abc_6362_n7911) );
	NAND2X1 NAND2X1_5353 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7911), .Y(dp.rf._abc_6362_n7912) );
	INVX1 INVX1_230 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<25>), .Y(dp.rf._abc_6362_n7913) );
	NOR2X1 NOR2X1_785 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7913), .Y(dp.rf._abc_6362_n7914) );
	NOR2X1 NOR2X1_786 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7912), .B(dp.rf._abc_6362_n7914), .Y(dp.rf._abc_6362_n7915) );
	NAND2X1 NAND2X1_5354 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<25>), .Y(dp.rf._abc_6362_n7916) );
	NAND2X1 NAND2X1_5355 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7916), .Y(dp.rf._abc_6362_n7917) );
	INVX1 INVX1_231 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<25>), .Y(dp.rf._abc_6362_n7918) );
	NOR2X1 NOR2X1_787 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n7918), .Y(dp.rf._abc_6362_n7919) );
	NOR2X1 NOR2X1_788 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7917), .B(dp.rf._abc_6362_n7919), .Y(dp.rf._abc_6362_n7920) );
	OR2X2 OR2X2_71 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7915), .B(dp.rf._abc_6362_n7920), .Y(dp.rf._abc_6362_n7921) );
	NAND2X1 NAND2X1_5356 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7921), .Y(dp.rf._abc_6362_n7922) );
	AND2X2 AND2X2_286 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7922), .B(instr[24]), .Y(dp.rf._abc_6362_n7923) );
	NAND2X1 NAND2X1_5357 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7910), .B(dp.rf._abc_6362_n7923), .Y(dp.rf._abc_6362_n7924) );
	NAND2X1 NAND2X1_5358 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7924), .Y(dp.rf._abc_6362_n7925) );
	NOR2X1 NOR2X1_789 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7898), .B(dp.rf._abc_6362_n7925), .Y(dp.rf._abc_6362_n7926) );
	NAND2X1 NAND2X1_5359 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<25>), .Y(dp.rf._abc_6362_n7927) );
	NAND2X1 NAND2X1_5360 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7928) );
	NAND2X1 NAND2X1_5361 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7927), .B(dp.rf._abc_6362_n7928), .Y(dp.rf._abc_6362_n7929) );
	NAND2X1 NAND2X1_5362 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7929), .Y(dp.rf._abc_6362_n7930) );
	NAND2X1 NAND2X1_5363 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<25>), .Y(dp.rf._abc_6362_n7931) );
	NAND2X1 NAND2X1_5364 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7932) );
	NAND2X1 NAND2X1_5365 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7931), .B(dp.rf._abc_6362_n7932), .Y(dp.rf._abc_6362_n7933) );
	NAND2X1 NAND2X1_5366 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7933), .Y(dp.rf._abc_6362_n7934) );
	AND2X2 AND2X2_287 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7930), .B(dp.rf._abc_6362_n7934), .Y(dp.rf._abc_6362_n7935) );
	NAND2X1 NAND2X1_5367 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n7935), .Y(dp.rf._abc_6362_n7936) );
	NAND2X1 NAND2X1_5368 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<25>), .Y(dp.rf._abc_6362_n7937) );
	NAND2X1 NAND2X1_5369 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7938) );
	NAND2X1 NAND2X1_5370 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7937), .B(dp.rf._abc_6362_n7938), .Y(dp.rf._abc_6362_n7939) );
	NAND2X1 NAND2X1_5371 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7939), .Y(dp.rf._abc_6362_n7940) );
	NAND2X1 NAND2X1_5372 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<25>), .Y(dp.rf._abc_6362_n7941) );
	NAND2X1 NAND2X1_5373 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7942) );
	NAND2X1 NAND2X1_5374 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7941), .B(dp.rf._abc_6362_n7942), .Y(dp.rf._abc_6362_n7943) );
	NAND2X1 NAND2X1_5375 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7943), .Y(dp.rf._abc_6362_n7944) );
	AND2X2 AND2X2_288 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7940), .B(dp.rf._abc_6362_n7944), .Y(dp.rf._abc_6362_n7945) );
	NAND2X1 NAND2X1_5376 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7945), .Y(dp.rf._abc_6362_n7946) );
	AND2X2 AND2X2_289 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7946), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n7947) );
	NAND2X1 NAND2X1_5377 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7936), .B(dp.rf._abc_6362_n7947), .Y(dp.rf._abc_6362_n7948) );
	NAND2X1 NAND2X1_5378 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7949) );
	NAND2X1 NAND2X1_5379 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<25>), .Y(dp.rf._abc_6362_n7950) );
	AND2X2 AND2X2_290 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7950), .B(instr[22]), .Y(dp.rf._abc_6362_n7951) );
	NAND2X1 NAND2X1_5380 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7949), .B(dp.rf._abc_6362_n7951), .Y(dp.rf._abc_6362_n7952) );
	NAND2X1 NAND2X1_5381 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7953) );
	NAND2X1 NAND2X1_5382 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<25>), .Y(dp.rf._abc_6362_n7954) );
	AND2X2 AND2X2_291 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7954), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7955) );
	NAND2X1 NAND2X1_5383 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7953), .B(dp.rf._abc_6362_n7955), .Y(dp.rf._abc_6362_n7956) );
	NAND2X1 NAND2X1_5384 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7952), .B(dp.rf._abc_6362_n7956), .Y(dp.rf._abc_6362_n7957) );
	AND2X2 AND2X2_292 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7957), .B(instr[23]), .Y(dp.rf._abc_6362_n7958) );
	NAND2X1 NAND2X1_5385 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7959) );
	NAND2X1 NAND2X1_5386 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<25>), .Y(dp.rf._abc_6362_n7960) );
	AND2X2 AND2X2_293 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7960), .B(instr[22]), .Y(dp.rf._abc_6362_n7961) );
	NAND2X1 NAND2X1_5387 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7959), .B(dp.rf._abc_6362_n7961), .Y(dp.rf._abc_6362_n7962) );
	NAND2X1 NAND2X1_5388 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<25>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7963) );
	NAND2X1 NAND2X1_5389 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<25>), .Y(dp.rf._abc_6362_n7964) );
	AND2X2 AND2X2_294 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7964), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n7965) );
	NAND2X1 NAND2X1_5390 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7963), .B(dp.rf._abc_6362_n7965), .Y(dp.rf._abc_6362_n7966) );
	NAND2X1 NAND2X1_5391 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7962), .B(dp.rf._abc_6362_n7966), .Y(dp.rf._abc_6362_n7967) );
	NAND2X1 NAND2X1_5392 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7967), .Y(dp.rf._abc_6362_n7968) );
	NAND2X1 NAND2X1_5393 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n7968), .Y(dp.rf._abc_6362_n7969) );
	NOR2X1 NOR2X1_790 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7958), .B(dp.rf._abc_6362_n7969), .Y(dp.rf._abc_6362_n7970) );
	NOR2X1 NOR2X1_791 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n7970), .Y(dp.rf._abc_6362_n7971) );
	NAND2X1 NAND2X1_5394 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7948), .B(dp.rf._abc_6362_n7971), .Y(dp.rf._abc_6362_n7972) );
	NAND2X1 NAND2X1_5395 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n7972), .Y(dp.rf._abc_6362_n7973) );
	NOR2X1 NOR2X1_792 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7926), .B(dp.rf._abc_6362_n7973), .Y(dp.srca_25_) );
	NAND2X1 NAND2X1_5396 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<26>), .Y(dp.rf._abc_6362_n7975) );
	NAND2X1 NAND2X1_5397 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7976) );
	NAND2X1 NAND2X1_5398 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7975), .B(dp.rf._abc_6362_n7976), .Y(dp.rf._abc_6362_n7977) );
	NAND2X1 NAND2X1_5399 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7977), .Y(dp.rf._abc_6362_n7978) );
	NAND2X1 NAND2X1_5400 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<26>), .Y(dp.rf._abc_6362_n7979) );
	NAND2X1 NAND2X1_5401 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7980) );
	NAND2X1 NAND2X1_5402 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7979), .B(dp.rf._abc_6362_n7980), .Y(dp.rf._abc_6362_n7981) );
	NAND2X1 NAND2X1_5403 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7981), .Y(dp.rf._abc_6362_n7982) );
	NAND2X1 NAND2X1_5404 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7978), .B(dp.rf._abc_6362_n7982), .Y(dp.rf._abc_6362_n7983) );
	NOR2X1 NOR2X1_793 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7983), .Y(dp.rf._abc_6362_n7984) );
	NAND2X1 NAND2X1_5405 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<26>), .Y(dp.rf._abc_6362_n7985) );
	NAND2X1 NAND2X1_5406 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7986) );
	NAND2X1 NAND2X1_5407 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7985), .B(dp.rf._abc_6362_n7986), .Y(dp.rf._abc_6362_n7987) );
	NAND2X1 NAND2X1_5408 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7987), .Y(dp.rf._abc_6362_n7988) );
	NAND2X1 NAND2X1_5409 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<26>), .Y(dp.rf._abc_6362_n7989) );
	NAND2X1 NAND2X1_5410 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7990) );
	NAND2X1 NAND2X1_5411 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7989), .B(dp.rf._abc_6362_n7990), .Y(dp.rf._abc_6362_n7991) );
	NAND2X1 NAND2X1_5412 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n7991), .Y(dp.rf._abc_6362_n7992) );
	AND2X2 AND2X2_295 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7988), .B(dp.rf._abc_6362_n7992), .Y(dp.rf._abc_6362_n7993) );
	NAND2X1 NAND2X1_5413 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n7993), .Y(dp.rf._abc_6362_n7994) );
	NAND2X1 NAND2X1_5414 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n7994), .Y(dp.rf._abc_6362_n7995) );
	NOR2X1 NOR2X1_794 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7984), .B(dp.rf._abc_6362_n7995), .Y(dp.rf._abc_6362_n7996) );
	NAND2X1 NAND2X1_5415 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<26>), .Y(dp.rf._abc_6362_n7997) );
	NAND2X1 NAND2X1_5416 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n7998) );
	NAND2X1 NAND2X1_5417 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7997), .B(dp.rf._abc_6362_n7998), .Y(dp.rf._abc_6362_n7999) );
	NAND2X1 NAND2X1_5418 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n7999), .Y(dp.rf._abc_6362_n8000) );
	NAND2X1 NAND2X1_5419 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<26>), .Y(dp.rf._abc_6362_n8001) );
	NAND2X1 NAND2X1_5420 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8002) );
	NAND2X1 NAND2X1_5421 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8001), .B(dp.rf._abc_6362_n8002), .Y(dp.rf._abc_6362_n8003) );
	NAND2X1 NAND2X1_5422 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8003), .Y(dp.rf._abc_6362_n8004) );
	NAND2X1 NAND2X1_5423 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8000), .B(dp.rf._abc_6362_n8004), .Y(dp.rf._abc_6362_n8005) );
	NAND2X1 NAND2X1_5424 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8005), .Y(dp.rf._abc_6362_n8006) );
	NAND2X1 NAND2X1_5425 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<26>), .Y(dp.rf._abc_6362_n8007) );
	NAND2X1 NAND2X1_5426 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8008) );
	NAND2X1 NAND2X1_5427 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8007), .B(dp.rf._abc_6362_n8008), .Y(dp.rf._abc_6362_n8009) );
	NAND2X1 NAND2X1_5428 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8009), .Y(dp.rf._abc_6362_n8010) );
	NAND2X1 NAND2X1_5429 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<26>), .Y(dp.rf._abc_6362_n8011) );
	NAND2X1 NAND2X1_5430 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8012) );
	NAND2X1 NAND2X1_5431 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8011), .B(dp.rf._abc_6362_n8012), .Y(dp.rf._abc_6362_n8013) );
	NAND2X1 NAND2X1_5432 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8013), .Y(dp.rf._abc_6362_n8014) );
	NAND2X1 NAND2X1_5433 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8010), .B(dp.rf._abc_6362_n8014), .Y(dp.rf._abc_6362_n8015) );
	NAND2X1 NAND2X1_5434 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8015), .Y(dp.rf._abc_6362_n8016) );
	NAND2X1 NAND2X1_5435 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8006), .B(dp.rf._abc_6362_n8016), .Y(dp.rf._abc_6362_n8017) );
	NAND2X1 NAND2X1_5436 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n8017), .Y(dp.rf._abc_6362_n8018) );
	NAND2X1 NAND2X1_5437 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n8018), .Y(dp.rf._abc_6362_n8019) );
	NOR2X1 NOR2X1_795 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n7996), .B(dp.rf._abc_6362_n8019), .Y(dp.rf._abc_6362_n8020) );
	NAND2X1 NAND2X1_5438 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<26>), .Y(dp.rf._abc_6362_n8021) );
	NAND2X1 NAND2X1_5439 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8022) );
	NAND2X1 NAND2X1_5440 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8021), .B(dp.rf._abc_6362_n8022), .Y(dp.rf._abc_6362_n8023) );
	NAND2X1 NAND2X1_5441 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8023), .Y(dp.rf._abc_6362_n8024) );
	NAND2X1 NAND2X1_5442 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<26>), .Y(dp.rf._abc_6362_n8025) );
	NAND2X1 NAND2X1_5443 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8026) );
	NAND2X1 NAND2X1_5444 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8025), .B(dp.rf._abc_6362_n8026), .Y(dp.rf._abc_6362_n8027) );
	NAND2X1 NAND2X1_5445 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8027), .Y(dp.rf._abc_6362_n8028) );
	NAND2X1 NAND2X1_5446 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8024), .B(dp.rf._abc_6362_n8028), .Y(dp.rf._abc_6362_n8029) );
	NAND2X1 NAND2X1_5447 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8029), .Y(dp.rf._abc_6362_n8030) );
	NAND2X1 NAND2X1_5448 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<26>), .Y(dp.rf._abc_6362_n8031) );
	NAND2X1 NAND2X1_5449 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8032) );
	NAND2X1 NAND2X1_5450 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8031), .B(dp.rf._abc_6362_n8032), .Y(dp.rf._abc_6362_n8033) );
	NAND2X1 NAND2X1_5451 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8033), .Y(dp.rf._abc_6362_n8034) );
	NAND2X1 NAND2X1_5452 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<26>), .Y(dp.rf._abc_6362_n8035) );
	NAND2X1 NAND2X1_5453 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8036) );
	NAND2X1 NAND2X1_5454 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8035), .B(dp.rf._abc_6362_n8036), .Y(dp.rf._abc_6362_n8037) );
	NAND2X1 NAND2X1_5455 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8037), .Y(dp.rf._abc_6362_n8038) );
	NAND2X1 NAND2X1_5456 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8034), .B(dp.rf._abc_6362_n8038), .Y(dp.rf._abc_6362_n8039) );
	NAND2X1 NAND2X1_5457 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8039), .Y(dp.rf._abc_6362_n8040) );
	NAND2X1 NAND2X1_5458 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8030), .B(dp.rf._abc_6362_n8040), .Y(dp.rf._abc_6362_n8041) );
	NAND2X1 NAND2X1_5459 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n8041), .Y(dp.rf._abc_6362_n8042) );
	NAND2X1 NAND2X1_5460 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8043) );
	NAND2X1 NAND2X1_5461 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<26>), .Y(dp.rf._abc_6362_n8044) );
	AND2X2 AND2X2_296 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8044), .B(instr[22]), .Y(dp.rf._abc_6362_n8045) );
	NAND2X1 NAND2X1_5462 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8043), .B(dp.rf._abc_6362_n8045), .Y(dp.rf._abc_6362_n8046) );
	NAND2X1 NAND2X1_5463 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8047) );
	NAND2X1 NAND2X1_5464 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<26>), .Y(dp.rf._abc_6362_n8048) );
	AND2X2 AND2X2_297 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8048), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8049) );
	NAND2X1 NAND2X1_5465 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8047), .B(dp.rf._abc_6362_n8049), .Y(dp.rf._abc_6362_n8050) );
	NAND2X1 NAND2X1_5466 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8046), .B(dp.rf._abc_6362_n8050), .Y(dp.rf._abc_6362_n8051) );
	AND2X2 AND2X2_298 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8051), .B(instr[23]), .Y(dp.rf._abc_6362_n8052) );
	NAND2X1 NAND2X1_5467 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8053) );
	NAND2X1 NAND2X1_5468 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<26>), .Y(dp.rf._abc_6362_n8054) );
	AND2X2 AND2X2_299 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8054), .B(instr[22]), .Y(dp.rf._abc_6362_n8055) );
	NAND2X1 NAND2X1_5469 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8053), .B(dp.rf._abc_6362_n8055), .Y(dp.rf._abc_6362_n8056) );
	NAND2X1 NAND2X1_5470 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<26>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8057) );
	NAND2X1 NAND2X1_5471 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<26>), .Y(dp.rf._abc_6362_n8058) );
	AND2X2 AND2X2_300 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8058), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8059) );
	NAND2X1 NAND2X1_5472 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8057), .B(dp.rf._abc_6362_n8059), .Y(dp.rf._abc_6362_n8060) );
	NAND2X1 NAND2X1_5473 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8056), .B(dp.rf._abc_6362_n8060), .Y(dp.rf._abc_6362_n8061) );
	NAND2X1 NAND2X1_5474 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8061), .Y(dp.rf._abc_6362_n8062) );
	NAND2X1 NAND2X1_5475 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n8062), .Y(dp.rf._abc_6362_n8063) );
	NOR2X1 NOR2X1_796 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8052), .B(dp.rf._abc_6362_n8063), .Y(dp.rf._abc_6362_n8064) );
	NOR2X1 NOR2X1_797 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n8064), .Y(dp.rf._abc_6362_n8065) );
	NAND2X1 NAND2X1_5476 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8042), .B(dp.rf._abc_6362_n8065), .Y(dp.rf._abc_6362_n8066) );
	NAND2X1 NAND2X1_5477 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n8066), .Y(dp.rf._abc_6362_n8067) );
	NOR2X1 NOR2X1_798 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8020), .B(dp.rf._abc_6362_n8067), .Y(dp.srca_26_) );
	NAND2X1 NAND2X1_5478 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<27>), .Y(dp.rf._abc_6362_n8069) );
	NAND2X1 NAND2X1_5479 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<27>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8070) );
	NAND2X1 NAND2X1_5480 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8069), .B(dp.rf._abc_6362_n8070), .Y(dp.rf._abc_6362_n8071) );
	NAND2X1 NAND2X1_5481 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8071), .Y(dp.rf._abc_6362_n8072) );
	NAND2X1 NAND2X1_5482 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<27>), .Y(dp.rf._abc_6362_n8073) );
	NAND2X1 NAND2X1_5483 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<27>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8074) );
	NAND2X1 NAND2X1_5484 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8073), .B(dp.rf._abc_6362_n8074), .Y(dp.rf._abc_6362_n8075) );
	NAND2X1 NAND2X1_5485 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8075), .Y(dp.rf._abc_6362_n8076) );
	NAND2X1 NAND2X1_5486 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8072), .B(dp.rf._abc_6362_n8076), .Y(dp.rf._abc_6362_n8077) );
	NOR2X1 NOR2X1_799 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8077), .Y(dp.rf._abc_6362_n8078) );
	NAND2X1 NAND2X1_5487 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<27>), .Y(dp.rf._abc_6362_n8079) );
	NAND2X1 NAND2X1_5488 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<27>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8080) );
	NAND2X1 NAND2X1_5489 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8079), .B(dp.rf._abc_6362_n8080), .Y(dp.rf._abc_6362_n8081) );
	NAND2X1 NAND2X1_5490 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8081), .Y(dp.rf._abc_6362_n8082) );
	NAND2X1 NAND2X1_5491 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<27>), .Y(dp.rf._abc_6362_n8083) );
	NAND2X1 NAND2X1_5492 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<27>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8084) );
	NAND2X1 NAND2X1_5493 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8083), .B(dp.rf._abc_6362_n8084), .Y(dp.rf._abc_6362_n8085) );
	NAND2X1 NAND2X1_5494 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8085), .Y(dp.rf._abc_6362_n8086) );
	AND2X2 AND2X2_301 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8082), .B(dp.rf._abc_6362_n8086), .Y(dp.rf._abc_6362_n8087) );
	NAND2X1 NAND2X1_5495 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8087), .Y(dp.rf._abc_6362_n8088) );
	NAND2X1 NAND2X1_5496 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n8088), .Y(dp.rf._abc_6362_n8089) );
	NOR2X1 NOR2X1_800 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8078), .B(dp.rf._abc_6362_n8089), .Y(dp.rf._abc_6362_n8090) );
	NAND2X1 NAND2X1_5497 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<27>), .Y(dp.rf._abc_6362_n8091) );
	NAND2X1 NAND2X1_5498 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<27>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8092) );
	NAND2X1 NAND2X1_5499 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8091), .B(dp.rf._abc_6362_n8092), .Y(dp.rf._abc_6362_n8093) );
	NAND2X1 NAND2X1_5500 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8093), .Y(dp.rf._abc_6362_n8094) );
	NAND2X1 NAND2X1_5501 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<27>), .Y(dp.rf._abc_6362_n8095) );
	NAND2X1 NAND2X1_5502 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<27>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8096) );
	NAND2X1 NAND2X1_5503 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8095), .B(dp.rf._abc_6362_n8096), .Y(dp.rf._abc_6362_n8097) );
	NAND2X1 NAND2X1_5504 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8097), .Y(dp.rf._abc_6362_n8098) );
	AND2X2 AND2X2_302 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8094), .B(dp.rf._abc_6362_n8098), .Y(dp.rf._abc_6362_n8099) );
	NAND2X1 NAND2X1_5505 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8099), .Y(dp.rf._abc_6362_n8100) );
	NAND2X1 NAND2X1_5506 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<27>), .Y(dp.rf._abc_6362_n8101) );
	NAND2X1 NAND2X1_5507 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8101), .Y(dp.rf._abc_6362_n8102) );
	AND2X2 AND2X2_303 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf.rf_2_<27>), .Y(dp.rf._abc_6362_n8103) );
	NOR2X1 NOR2X1_801 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8102), .B(dp.rf._abc_6362_n8103), .Y(dp.rf._abc_6362_n8104) );
	NAND2X1 NAND2X1_5508 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<27>), .Y(dp.rf._abc_6362_n8105) );
	NAND2X1 NAND2X1_5509 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8105), .Y(dp.rf._abc_6362_n8106) );
	INVX1 INVX1_232 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<27>), .Y(dp.rf._abc_6362_n8107) );
	NOR2X1 NOR2X1_802 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8107), .Y(dp.rf._abc_6362_n8108) );
	NOR2X1 NOR2X1_803 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8106), .B(dp.rf._abc_6362_n8108), .Y(dp.rf._abc_6362_n8109) );
	OR2X2 OR2X2_72 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8104), .B(dp.rf._abc_6362_n8109), .Y(dp.rf._abc_6362_n8110) );
	NAND2X1 NAND2X1_5510 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8110), .Y(dp.rf._abc_6362_n8111) );
	AND2X2 AND2X2_304 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8111), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n8112) );
	NAND2X1 NAND2X1_5511 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8100), .B(dp.rf._abc_6362_n8112), .Y(dp.rf._abc_6362_n8113) );
	NAND2X1 NAND2X1_5512 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n8113), .Y(dp.rf._abc_6362_n8114) );
	NOR2X1 NOR2X1_804 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8090), .B(dp.rf._abc_6362_n8114), .Y(dp.rf._abc_6362_n8115) );
	NAND2X1 NAND2X1_5513 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<27>), .Y(dp.rf._abc_6362_n8116) );
	NAND2X1 NAND2X1_5514 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8116), .Y(dp.rf._abc_6362_n8117) );
	INVX1 INVX1_233 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<27>), .Y(dp.rf._abc_6362_n8118) );
	NOR2X1 NOR2X1_805 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8118), .Y(dp.rf._abc_6362_n8119) );
	NOR2X1 NOR2X1_806 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8117), .B(dp.rf._abc_6362_n8119), .Y(dp.rf._abc_6362_n8120) );
	NAND2X1 NAND2X1_5515 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<27>), .Y(dp.rf._abc_6362_n8121) );
	NAND2X1 NAND2X1_5516 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8121), .Y(dp.rf._abc_6362_n8122) );
	INVX1 INVX1_234 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<27>), .Y(dp.rf._abc_6362_n8123) );
	NOR2X1 NOR2X1_807 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8123), .Y(dp.rf._abc_6362_n8124) );
	NOR2X1 NOR2X1_808 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8122), .B(dp.rf._abc_6362_n8124), .Y(dp.rf._abc_6362_n8125) );
	OR2X2 OR2X2_73 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8120), .B(dp.rf._abc_6362_n8125), .Y(dp.rf._abc_6362_n8126) );
	NAND2X1 NAND2X1_5517 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8126), .Y(dp.rf._abc_6362_n8127) );
	NAND2X1 NAND2X1_5518 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<27>), .Y(dp.rf._abc_6362_n8128) );
	NAND2X1 NAND2X1_5519 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8128), .Y(dp.rf._abc_6362_n8129) );
	INVX1 INVX1_235 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<27>), .Y(dp.rf._abc_6362_n8130) );
	NOR2X1 NOR2X1_809 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8130), .Y(dp.rf._abc_6362_n8131) );
	NOR2X1 NOR2X1_810 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8129), .B(dp.rf._abc_6362_n8131), .Y(dp.rf._abc_6362_n8132) );
	NAND2X1 NAND2X1_5520 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<27>), .Y(dp.rf._abc_6362_n8133) );
	NAND2X1 NAND2X1_5521 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8133), .Y(dp.rf._abc_6362_n8134) );
	INVX1 INVX1_236 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<27>), .Y(dp.rf._abc_6362_n8135) );
	NOR2X1 NOR2X1_811 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8135), .Y(dp.rf._abc_6362_n8136) );
	NOR2X1 NOR2X1_812 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8134), .B(dp.rf._abc_6362_n8136), .Y(dp.rf._abc_6362_n8137) );
	OR2X2 OR2X2_74 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8132), .B(dp.rf._abc_6362_n8137), .Y(dp.rf._abc_6362_n8138) );
	NAND2X1 NAND2X1_5522 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8138), .Y(dp.rf._abc_6362_n8139) );
	AND2X2 AND2X2_305 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8139), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n8140) );
	NAND2X1 NAND2X1_5523 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8127), .B(dp.rf._abc_6362_n8140), .Y(dp.rf._abc_6362_n8141) );
	NAND2X1 NAND2X1_5524 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<27>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8142) );
	NAND2X1 NAND2X1_5525 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<27>), .Y(dp.rf._abc_6362_n8143) );
	AND2X2 AND2X2_306 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8143), .B(instr[22]), .Y(dp.rf._abc_6362_n8144) );
	NAND2X1 NAND2X1_5526 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8142), .B(dp.rf._abc_6362_n8144), .Y(dp.rf._abc_6362_n8145) );
	NAND2X1 NAND2X1_5527 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<27>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8146) );
	NAND2X1 NAND2X1_5528 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<27>), .Y(dp.rf._abc_6362_n8147) );
	AND2X2 AND2X2_307 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8147), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8148) );
	NAND2X1 NAND2X1_5529 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8146), .B(dp.rf._abc_6362_n8148), .Y(dp.rf._abc_6362_n8149) );
	NAND2X1 NAND2X1_5530 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8145), .B(dp.rf._abc_6362_n8149), .Y(dp.rf._abc_6362_n8150) );
	AND2X2 AND2X2_308 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8150), .B(instr[23]), .Y(dp.rf._abc_6362_n8151) );
	NAND2X1 NAND2X1_5531 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<27>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8152) );
	NAND2X1 NAND2X1_5532 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<27>), .Y(dp.rf._abc_6362_n8153) );
	AND2X2 AND2X2_309 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8153), .B(instr[22]), .Y(dp.rf._abc_6362_n8154) );
	NAND2X1 NAND2X1_5533 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8152), .B(dp.rf._abc_6362_n8154), .Y(dp.rf._abc_6362_n8155) );
	NAND2X1 NAND2X1_5534 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<27>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8156) );
	NAND2X1 NAND2X1_5535 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<27>), .Y(dp.rf._abc_6362_n8157) );
	AND2X2 AND2X2_310 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8157), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8158) );
	NAND2X1 NAND2X1_5536 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8156), .B(dp.rf._abc_6362_n8158), .Y(dp.rf._abc_6362_n8159) );
	NAND2X1 NAND2X1_5537 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8155), .B(dp.rf._abc_6362_n8159), .Y(dp.rf._abc_6362_n8160) );
	NAND2X1 NAND2X1_5538 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8160), .Y(dp.rf._abc_6362_n8161) );
	NAND2X1 NAND2X1_5539 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n8161), .Y(dp.rf._abc_6362_n8162) );
	NOR2X1 NOR2X1_813 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8151), .B(dp.rf._abc_6362_n8162), .Y(dp.rf._abc_6362_n8163) );
	NOR2X1 NOR2X1_814 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n8163), .Y(dp.rf._abc_6362_n8164) );
	NAND2X1 NAND2X1_5540 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8141), .B(dp.rf._abc_6362_n8164), .Y(dp.rf._abc_6362_n8165) );
	NAND2X1 NAND2X1_5541 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n8165), .Y(dp.rf._abc_6362_n8166) );
	NOR2X1 NOR2X1_815 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8115), .B(dp.rf._abc_6362_n8166), .Y(dp.srca_27_) );
	NAND2X1 NAND2X1_5542 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<28>), .Y(dp.rf._abc_6362_n8168) );
	NAND2X1 NAND2X1_5543 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8169) );
	NAND2X1 NAND2X1_5544 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8168), .B(dp.rf._abc_6362_n8169), .Y(dp.rf._abc_6362_n8170) );
	NAND2X1 NAND2X1_5545 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8170), .Y(dp.rf._abc_6362_n8171) );
	NAND2X1 NAND2X1_5546 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<28>), .Y(dp.rf._abc_6362_n8172) );
	NAND2X1 NAND2X1_5547 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8173) );
	NAND2X1 NAND2X1_5548 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8172), .B(dp.rf._abc_6362_n8173), .Y(dp.rf._abc_6362_n8174) );
	NAND2X1 NAND2X1_5549 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8174), .Y(dp.rf._abc_6362_n8175) );
	NAND2X1 NAND2X1_5550 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8171), .B(dp.rf._abc_6362_n8175), .Y(dp.rf._abc_6362_n8176) );
	NOR2X1 NOR2X1_816 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8176), .Y(dp.rf._abc_6362_n8177) );
	NAND2X1 NAND2X1_5551 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<28>), .Y(dp.rf._abc_6362_n8178) );
	NAND2X1 NAND2X1_5552 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8179) );
	NAND2X1 NAND2X1_5553 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8178), .B(dp.rf._abc_6362_n8179), .Y(dp.rf._abc_6362_n8180) );
	NAND2X1 NAND2X1_5554 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8180), .Y(dp.rf._abc_6362_n8181) );
	NAND2X1 NAND2X1_5555 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<28>), .Y(dp.rf._abc_6362_n8182) );
	NAND2X1 NAND2X1_5556 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8183) );
	NAND2X1 NAND2X1_5557 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8182), .B(dp.rf._abc_6362_n8183), .Y(dp.rf._abc_6362_n8184) );
	NAND2X1 NAND2X1_5558 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8184), .Y(dp.rf._abc_6362_n8185) );
	AND2X2 AND2X2_311 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8181), .B(dp.rf._abc_6362_n8185), .Y(dp.rf._abc_6362_n8186) );
	NAND2X1 NAND2X1_5559 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8186), .Y(dp.rf._abc_6362_n8187) );
	NAND2X1 NAND2X1_5560 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n8187), .Y(dp.rf._abc_6362_n8188) );
	NOR2X1 NOR2X1_817 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8177), .B(dp.rf._abc_6362_n8188), .Y(dp.rf._abc_6362_n8189) );
	NAND2X1 NAND2X1_5561 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<28>), .Y(dp.rf._abc_6362_n8190) );
	NAND2X1 NAND2X1_5562 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8191) );
	NAND2X1 NAND2X1_5563 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8190), .B(dp.rf._abc_6362_n8191), .Y(dp.rf._abc_6362_n8192) );
	NAND2X1 NAND2X1_5564 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8192), .Y(dp.rf._abc_6362_n8193) );
	NAND2X1 NAND2X1_5565 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<28>), .Y(dp.rf._abc_6362_n8194) );
	NAND2X1 NAND2X1_5566 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8195) );
	NAND2X1 NAND2X1_5567 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8194), .B(dp.rf._abc_6362_n8195), .Y(dp.rf._abc_6362_n8196) );
	NAND2X1 NAND2X1_5568 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8196), .Y(dp.rf._abc_6362_n8197) );
	NAND2X1 NAND2X1_5569 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8193), .B(dp.rf._abc_6362_n8197), .Y(dp.rf._abc_6362_n8198) );
	NAND2X1 NAND2X1_5570 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8198), .Y(dp.rf._abc_6362_n8199) );
	NAND2X1 NAND2X1_5571 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<28>), .Y(dp.rf._abc_6362_n8200) );
	NAND2X1 NAND2X1_5572 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8201) );
	NAND2X1 NAND2X1_5573 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8200), .B(dp.rf._abc_6362_n8201), .Y(dp.rf._abc_6362_n8202) );
	NAND2X1 NAND2X1_5574 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8202), .Y(dp.rf._abc_6362_n8203) );
	NAND2X1 NAND2X1_5575 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<28>), .Y(dp.rf._abc_6362_n8204) );
	NAND2X1 NAND2X1_5576 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8205) );
	NAND2X1 NAND2X1_5577 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8204), .B(dp.rf._abc_6362_n8205), .Y(dp.rf._abc_6362_n8206) );
	NAND2X1 NAND2X1_5578 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8206), .Y(dp.rf._abc_6362_n8207) );
	NAND2X1 NAND2X1_5579 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8203), .B(dp.rf._abc_6362_n8207), .Y(dp.rf._abc_6362_n8208) );
	NAND2X1 NAND2X1_5580 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8208), .Y(dp.rf._abc_6362_n8209) );
	NAND2X1 NAND2X1_5581 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8199), .B(dp.rf._abc_6362_n8209), .Y(dp.rf._abc_6362_n8210) );
	NAND2X1 NAND2X1_5582 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n8210), .Y(dp.rf._abc_6362_n8211) );
	NAND2X1 NAND2X1_5583 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n8211), .Y(dp.rf._abc_6362_n8212) );
	NOR2X1 NOR2X1_818 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8189), .B(dp.rf._abc_6362_n8212), .Y(dp.rf._abc_6362_n8213) );
	NAND2X1 NAND2X1_5584 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<28>), .Y(dp.rf._abc_6362_n8214) );
	NAND2X1 NAND2X1_5585 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8214), .Y(dp.rf._abc_6362_n8215) );
	INVX1 INVX1_237 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<28>), .Y(dp.rf._abc_6362_n8216) );
	NOR2X1 NOR2X1_819 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8216), .Y(dp.rf._abc_6362_n8217) );
	NOR2X1 NOR2X1_820 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8215), .B(dp.rf._abc_6362_n8217), .Y(dp.rf._abc_6362_n8218) );
	NAND2X1 NAND2X1_5586 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<28>), .Y(dp.rf._abc_6362_n8219) );
	NAND2X1 NAND2X1_5587 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8219), .Y(dp.rf._abc_6362_n8220) );
	INVX1 INVX1_238 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<28>), .Y(dp.rf._abc_6362_n8221) );
	NOR2X1 NOR2X1_821 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8221), .Y(dp.rf._abc_6362_n8222) );
	NOR2X1 NOR2X1_822 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8220), .B(dp.rf._abc_6362_n8222), .Y(dp.rf._abc_6362_n8223) );
	OR2X2 OR2X2_75 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8218), .B(dp.rf._abc_6362_n8223), .Y(dp.rf._abc_6362_n8224) );
	NAND2X1 NAND2X1_5588 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8224), .Y(dp.rf._abc_6362_n8225) );
	NAND2X1 NAND2X1_5589 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<28>), .Y(dp.rf._abc_6362_n8226) );
	NAND2X1 NAND2X1_5590 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8226), .Y(dp.rf._abc_6362_n8227) );
	INVX1 INVX1_239 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<28>), .Y(dp.rf._abc_6362_n8228) );
	NOR2X1 NOR2X1_823 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8228), .Y(dp.rf._abc_6362_n8229) );
	NOR2X1 NOR2X1_824 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8227), .B(dp.rf._abc_6362_n8229), .Y(dp.rf._abc_6362_n8230) );
	NAND2X1 NAND2X1_5591 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<28>), .Y(dp.rf._abc_6362_n8231) );
	NAND2X1 NAND2X1_5592 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8231), .Y(dp.rf._abc_6362_n8232) );
	INVX1 INVX1_240 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<28>), .Y(dp.rf._abc_6362_n8233) );
	NOR2X1 NOR2X1_825 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8233), .Y(dp.rf._abc_6362_n8234) );
	NOR2X1 NOR2X1_826 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8232), .B(dp.rf._abc_6362_n8234), .Y(dp.rf._abc_6362_n8235) );
	OR2X2 OR2X2_76 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8230), .B(dp.rf._abc_6362_n8235), .Y(dp.rf._abc_6362_n8236) );
	NAND2X1 NAND2X1_5593 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8236), .Y(dp.rf._abc_6362_n8237) );
	AND2X2 AND2X2_312 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8237), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n8238) );
	NAND2X1 NAND2X1_5594 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8225), .B(dp.rf._abc_6362_n8238), .Y(dp.rf._abc_6362_n8239) );
	NAND2X1 NAND2X1_5595 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8240) );
	NAND2X1 NAND2X1_5596 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<28>), .Y(dp.rf._abc_6362_n8241) );
	AND2X2 AND2X2_313 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8241), .B(instr[22]), .Y(dp.rf._abc_6362_n8242) );
	NAND2X1 NAND2X1_5597 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8240), .B(dp.rf._abc_6362_n8242), .Y(dp.rf._abc_6362_n8243) );
	NAND2X1 NAND2X1_5598 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8244) );
	NAND2X1 NAND2X1_5599 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<28>), .Y(dp.rf._abc_6362_n8245) );
	AND2X2 AND2X2_314 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8245), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8246) );
	NAND2X1 NAND2X1_5600 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8244), .B(dp.rf._abc_6362_n8246), .Y(dp.rf._abc_6362_n8247) );
	NAND2X1 NAND2X1_5601 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8243), .B(dp.rf._abc_6362_n8247), .Y(dp.rf._abc_6362_n8248) );
	AND2X2 AND2X2_315 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8248), .B(instr[23]), .Y(dp.rf._abc_6362_n8249) );
	NAND2X1 NAND2X1_5602 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8250) );
	NAND2X1 NAND2X1_5603 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<28>), .Y(dp.rf._abc_6362_n8251) );
	AND2X2 AND2X2_316 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8251), .B(instr[22]), .Y(dp.rf._abc_6362_n8252) );
	NAND2X1 NAND2X1_5604 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8250), .B(dp.rf._abc_6362_n8252), .Y(dp.rf._abc_6362_n8253) );
	NAND2X1 NAND2X1_5605 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<28>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8254) );
	NAND2X1 NAND2X1_5606 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<28>), .Y(dp.rf._abc_6362_n8255) );
	AND2X2 AND2X2_317 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8255), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8256) );
	NAND2X1 NAND2X1_5607 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8254), .B(dp.rf._abc_6362_n8256), .Y(dp.rf._abc_6362_n8257) );
	NAND2X1 NAND2X1_5608 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8253), .B(dp.rf._abc_6362_n8257), .Y(dp.rf._abc_6362_n8258) );
	NAND2X1 NAND2X1_5609 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8258), .Y(dp.rf._abc_6362_n8259) );
	NAND2X1 NAND2X1_5610 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n8259), .Y(dp.rf._abc_6362_n8260) );
	NOR2X1 NOR2X1_827 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8249), .B(dp.rf._abc_6362_n8260), .Y(dp.rf._abc_6362_n8261) );
	NOR2X1 NOR2X1_828 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n8261), .Y(dp.rf._abc_6362_n8262) );
	NAND2X1 NAND2X1_5611 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8239), .B(dp.rf._abc_6362_n8262), .Y(dp.rf._abc_6362_n8263) );
	NAND2X1 NAND2X1_5612 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n8263), .Y(dp.rf._abc_6362_n8264) );
	NOR2X1 NOR2X1_829 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8213), .B(dp.rf._abc_6362_n8264), .Y(dp.srca_28_) );
	NAND2X1 NAND2X1_5613 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<29>), .Y(dp.rf._abc_6362_n8266) );
	NAND2X1 NAND2X1_5614 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<29>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8267) );
	NAND2X1 NAND2X1_5615 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8266), .B(dp.rf._abc_6362_n8267), .Y(dp.rf._abc_6362_n8268) );
	NAND2X1 NAND2X1_5616 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8268), .Y(dp.rf._abc_6362_n8269) );
	NAND2X1 NAND2X1_5617 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<29>), .Y(dp.rf._abc_6362_n8270) );
	NAND2X1 NAND2X1_5618 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<29>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8271) );
	NAND2X1 NAND2X1_5619 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8270), .B(dp.rf._abc_6362_n8271), .Y(dp.rf._abc_6362_n8272) );
	NAND2X1 NAND2X1_5620 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8272), .Y(dp.rf._abc_6362_n8273) );
	NAND2X1 NAND2X1_5621 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8269), .B(dp.rf._abc_6362_n8273), .Y(dp.rf._abc_6362_n8274) );
	NOR2X1 NOR2X1_830 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8274), .Y(dp.rf._abc_6362_n8275) );
	NAND2X1 NAND2X1_5622 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<29>), .Y(dp.rf._abc_6362_n8276) );
	NAND2X1 NAND2X1_5623 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<29>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8277) );
	NAND2X1 NAND2X1_5624 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8276), .B(dp.rf._abc_6362_n8277), .Y(dp.rf._abc_6362_n8278) );
	NAND2X1 NAND2X1_5625 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8278), .Y(dp.rf._abc_6362_n8279) );
	NAND2X1 NAND2X1_5626 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<29>), .Y(dp.rf._abc_6362_n8280) );
	NAND2X1 NAND2X1_5627 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<29>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8281) );
	NAND2X1 NAND2X1_5628 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8280), .B(dp.rf._abc_6362_n8281), .Y(dp.rf._abc_6362_n8282) );
	NAND2X1 NAND2X1_5629 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8282), .Y(dp.rf._abc_6362_n8283) );
	AND2X2 AND2X2_318 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8279), .B(dp.rf._abc_6362_n8283), .Y(dp.rf._abc_6362_n8284) );
	NAND2X1 NAND2X1_5630 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8284), .Y(dp.rf._abc_6362_n8285) );
	NAND2X1 NAND2X1_5631 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n8285), .Y(dp.rf._abc_6362_n8286) );
	NOR2X1 NOR2X1_831 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8275), .B(dp.rf._abc_6362_n8286), .Y(dp.rf._abc_6362_n8287) );
	NAND2X1 NAND2X1_5632 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<29>), .Y(dp.rf._abc_6362_n8288) );
	NAND2X1 NAND2X1_5633 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<29>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8289) );
	NAND2X1 NAND2X1_5634 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8288), .B(dp.rf._abc_6362_n8289), .Y(dp.rf._abc_6362_n8290) );
	NAND2X1 NAND2X1_5635 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8290), .Y(dp.rf._abc_6362_n8291) );
	NAND2X1 NAND2X1_5636 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<29>), .Y(dp.rf._abc_6362_n8292) );
	NAND2X1 NAND2X1_5637 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<29>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8293) );
	NAND2X1 NAND2X1_5638 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8292), .B(dp.rf._abc_6362_n8293), .Y(dp.rf._abc_6362_n8294) );
	NAND2X1 NAND2X1_5639 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8294), .Y(dp.rf._abc_6362_n8295) );
	AND2X2 AND2X2_319 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8291), .B(dp.rf._abc_6362_n8295), .Y(dp.rf._abc_6362_n8296) );
	NAND2X1 NAND2X1_5640 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8296), .Y(dp.rf._abc_6362_n8297) );
	NAND2X1 NAND2X1_5641 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<29>), .Y(dp.rf._abc_6362_n8298) );
	NAND2X1 NAND2X1_5642 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8298), .Y(dp.rf._abc_6362_n8299) );
	AND2X2 AND2X2_320 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5338), .B(dp.rf.rf_2_<29>), .Y(dp.rf._abc_6362_n8300) );
	NOR2X1 NOR2X1_832 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8299), .B(dp.rf._abc_6362_n8300), .Y(dp.rf._abc_6362_n8301) );
	NAND2X1 NAND2X1_5643 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<29>), .Y(dp.rf._abc_6362_n8302) );
	NAND2X1 NAND2X1_5644 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8302), .Y(dp.rf._abc_6362_n8303) );
	INVX1 INVX1_241 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<29>), .Y(dp.rf._abc_6362_n8304) );
	NOR2X1 NOR2X1_833 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8304), .Y(dp.rf._abc_6362_n8305) );
	NOR2X1 NOR2X1_834 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8303), .B(dp.rf._abc_6362_n8305), .Y(dp.rf._abc_6362_n8306) );
	OR2X2 OR2X2_77 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8301), .B(dp.rf._abc_6362_n8306), .Y(dp.rf._abc_6362_n8307) );
	NAND2X1 NAND2X1_5645 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8307), .Y(dp.rf._abc_6362_n8308) );
	AND2X2 AND2X2_321 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8308), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n8309) );
	NAND2X1 NAND2X1_5646 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8297), .B(dp.rf._abc_6362_n8309), .Y(dp.rf._abc_6362_n8310) );
	NAND2X1 NAND2X1_5647 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n8310), .Y(dp.rf._abc_6362_n8311) );
	NOR2X1 NOR2X1_835 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8287), .B(dp.rf._abc_6362_n8311), .Y(dp.rf._abc_6362_n8312) );
	NAND2X1 NAND2X1_5648 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<29>), .Y(dp.rf._abc_6362_n8313) );
	NAND2X1 NAND2X1_5649 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8313), .Y(dp.rf._abc_6362_n8314) );
	INVX1 INVX1_242 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<29>), .Y(dp.rf._abc_6362_n8315) );
	NOR2X1 NOR2X1_836 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8315), .Y(dp.rf._abc_6362_n8316) );
	NOR2X1 NOR2X1_837 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8314), .B(dp.rf._abc_6362_n8316), .Y(dp.rf._abc_6362_n8317) );
	NAND2X1 NAND2X1_5650 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<29>), .Y(dp.rf._abc_6362_n8318) );
	NAND2X1 NAND2X1_5651 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8318), .Y(dp.rf._abc_6362_n8319) );
	INVX1 INVX1_243 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<29>), .Y(dp.rf._abc_6362_n8320) );
	NOR2X1 NOR2X1_838 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8320), .Y(dp.rf._abc_6362_n8321) );
	NOR2X1 NOR2X1_839 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8319), .B(dp.rf._abc_6362_n8321), .Y(dp.rf._abc_6362_n8322) );
	OR2X2 OR2X2_78 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8317), .B(dp.rf._abc_6362_n8322), .Y(dp.rf._abc_6362_n8323) );
	NAND2X1 NAND2X1_5652 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8323), .Y(dp.rf._abc_6362_n8324) );
	NAND2X1 NAND2X1_5653 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<29>), .Y(dp.rf._abc_6362_n8325) );
	NAND2X1 NAND2X1_5654 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8325), .Y(dp.rf._abc_6362_n8326) );
	INVX1 INVX1_244 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<29>), .Y(dp.rf._abc_6362_n8327) );
	NOR2X1 NOR2X1_840 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8327), .Y(dp.rf._abc_6362_n8328) );
	NOR2X1 NOR2X1_841 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8326), .B(dp.rf._abc_6362_n8328), .Y(dp.rf._abc_6362_n8329) );
	NAND2X1 NAND2X1_5655 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<29>), .Y(dp.rf._abc_6362_n8330) );
	NAND2X1 NAND2X1_5656 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8330), .Y(dp.rf._abc_6362_n8331) );
	INVX1 INVX1_245 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<29>), .Y(dp.rf._abc_6362_n8332) );
	NOR2X1 NOR2X1_842 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8332), .Y(dp.rf._abc_6362_n8333) );
	NOR2X1 NOR2X1_843 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8331), .B(dp.rf._abc_6362_n8333), .Y(dp.rf._abc_6362_n8334) );
	OR2X2 OR2X2_79 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8329), .B(dp.rf._abc_6362_n8334), .Y(dp.rf._abc_6362_n8335) );
	NAND2X1 NAND2X1_5657 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8335), .Y(dp.rf._abc_6362_n8336) );
	AND2X2 AND2X2_322 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8336), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n8337) );
	NAND2X1 NAND2X1_5658 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8324), .B(dp.rf._abc_6362_n8337), .Y(dp.rf._abc_6362_n8338) );
	NAND2X1 NAND2X1_5659 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<29>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8339) );
	NAND2X1 NAND2X1_5660 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<29>), .Y(dp.rf._abc_6362_n8340) );
	AND2X2 AND2X2_323 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8340), .B(instr[22]), .Y(dp.rf._abc_6362_n8341) );
	NAND2X1 NAND2X1_5661 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8339), .B(dp.rf._abc_6362_n8341), .Y(dp.rf._abc_6362_n8342) );
	NAND2X1 NAND2X1_5662 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<29>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8343) );
	NAND2X1 NAND2X1_5663 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<29>), .Y(dp.rf._abc_6362_n8344) );
	AND2X2 AND2X2_324 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8344), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8345) );
	NAND2X1 NAND2X1_5664 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8343), .B(dp.rf._abc_6362_n8345), .Y(dp.rf._abc_6362_n8346) );
	NAND2X1 NAND2X1_5665 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8342), .B(dp.rf._abc_6362_n8346), .Y(dp.rf._abc_6362_n8347) );
	AND2X2 AND2X2_325 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8347), .B(instr[23]), .Y(dp.rf._abc_6362_n8348) );
	NAND2X1 NAND2X1_5666 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<29>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8349) );
	NAND2X1 NAND2X1_5667 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<29>), .Y(dp.rf._abc_6362_n8350) );
	AND2X2 AND2X2_326 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8350), .B(instr[22]), .Y(dp.rf._abc_6362_n8351) );
	NAND2X1 NAND2X1_5668 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8349), .B(dp.rf._abc_6362_n8351), .Y(dp.rf._abc_6362_n8352) );
	NAND2X1 NAND2X1_5669 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<29>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8353) );
	NAND2X1 NAND2X1_5670 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<29>), .Y(dp.rf._abc_6362_n8354) );
	AND2X2 AND2X2_327 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8354), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8355) );
	NAND2X1 NAND2X1_5671 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8353), .B(dp.rf._abc_6362_n8355), .Y(dp.rf._abc_6362_n8356) );
	NAND2X1 NAND2X1_5672 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8352), .B(dp.rf._abc_6362_n8356), .Y(dp.rf._abc_6362_n8357) );
	NAND2X1 NAND2X1_5673 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8357), .Y(dp.rf._abc_6362_n8358) );
	NAND2X1 NAND2X1_5674 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n8358), .Y(dp.rf._abc_6362_n8359) );
	NOR2X1 NOR2X1_844 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8348), .B(dp.rf._abc_6362_n8359), .Y(dp.rf._abc_6362_n8360) );
	NOR2X1 NOR2X1_845 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n8360), .Y(dp.rf._abc_6362_n8361) );
	NAND2X1 NAND2X1_5675 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8338), .B(dp.rf._abc_6362_n8361), .Y(dp.rf._abc_6362_n8362) );
	NAND2X1 NAND2X1_5676 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n8362), .Y(dp.rf._abc_6362_n8363) );
	NOR2X1 NOR2X1_846 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8312), .B(dp.rf._abc_6362_n8363), .Y(dp.srca_29_) );
	NAND2X1 NAND2X1_5677 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<30>), .Y(dp.rf._abc_6362_n8365) );
	NAND2X1 NAND2X1_5678 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8366) );
	NAND2X1 NAND2X1_5679 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8365), .B(dp.rf._abc_6362_n8366), .Y(dp.rf._abc_6362_n8367) );
	NAND2X1 NAND2X1_5680 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8367), .Y(dp.rf._abc_6362_n8368) );
	NAND2X1 NAND2X1_5681 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<30>), .Y(dp.rf._abc_6362_n8369) );
	NAND2X1 NAND2X1_5682 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8370) );
	NAND2X1 NAND2X1_5683 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8369), .B(dp.rf._abc_6362_n8370), .Y(dp.rf._abc_6362_n8371) );
	NAND2X1 NAND2X1_5684 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8371), .Y(dp.rf._abc_6362_n8372) );
	NAND2X1 NAND2X1_5685 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8368), .B(dp.rf._abc_6362_n8372), .Y(dp.rf._abc_6362_n8373) );
	NOR2X1 NOR2X1_847 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8373), .Y(dp.rf._abc_6362_n8374) );
	NAND2X1 NAND2X1_5686 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<30>), .Y(dp.rf._abc_6362_n8375) );
	NAND2X1 NAND2X1_5687 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8376) );
	NAND2X1 NAND2X1_5688 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8375), .B(dp.rf._abc_6362_n8376), .Y(dp.rf._abc_6362_n8377) );
	NAND2X1 NAND2X1_5689 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8377), .Y(dp.rf._abc_6362_n8378) );
	NAND2X1 NAND2X1_5690 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<30>), .Y(dp.rf._abc_6362_n8379) );
	NAND2X1 NAND2X1_5691 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8380) );
	NAND2X1 NAND2X1_5692 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8379), .B(dp.rf._abc_6362_n8380), .Y(dp.rf._abc_6362_n8381) );
	NAND2X1 NAND2X1_5693 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8381), .Y(dp.rf._abc_6362_n8382) );
	AND2X2 AND2X2_328 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8378), .B(dp.rf._abc_6362_n8382), .Y(dp.rf._abc_6362_n8383) );
	NAND2X1 NAND2X1_5694 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8383), .Y(dp.rf._abc_6362_n8384) );
	NAND2X1 NAND2X1_5695 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n8384), .Y(dp.rf._abc_6362_n8385) );
	NOR2X1 NOR2X1_848 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8374), .B(dp.rf._abc_6362_n8385), .Y(dp.rf._abc_6362_n8386) );
	NAND2X1 NAND2X1_5696 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<30>), .Y(dp.rf._abc_6362_n8387) );
	NAND2X1 NAND2X1_5697 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8388) );
	NAND2X1 NAND2X1_5698 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8387), .B(dp.rf._abc_6362_n8388), .Y(dp.rf._abc_6362_n8389) );
	NAND2X1 NAND2X1_5699 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8389), .Y(dp.rf._abc_6362_n8390) );
	NAND2X1 NAND2X1_5700 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<30>), .Y(dp.rf._abc_6362_n8391) );
	NAND2X1 NAND2X1_5701 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8392) );
	NAND2X1 NAND2X1_5702 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8391), .B(dp.rf._abc_6362_n8392), .Y(dp.rf._abc_6362_n8393) );
	NAND2X1 NAND2X1_5703 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8393), .Y(dp.rf._abc_6362_n8394) );
	NAND2X1 NAND2X1_5704 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8390), .B(dp.rf._abc_6362_n8394), .Y(dp.rf._abc_6362_n8395) );
	NAND2X1 NAND2X1_5705 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8395), .Y(dp.rf._abc_6362_n8396) );
	NAND2X1 NAND2X1_5706 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<30>), .Y(dp.rf._abc_6362_n8397) );
	NAND2X1 NAND2X1_5707 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8398) );
	NAND2X1 NAND2X1_5708 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8397), .B(dp.rf._abc_6362_n8398), .Y(dp.rf._abc_6362_n8399) );
	NAND2X1 NAND2X1_5709 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8399), .Y(dp.rf._abc_6362_n8400) );
	NAND2X1 NAND2X1_5710 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<30>), .Y(dp.rf._abc_6362_n8401) );
	NAND2X1 NAND2X1_5711 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8402) );
	NAND2X1 NAND2X1_5712 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8401), .B(dp.rf._abc_6362_n8402), .Y(dp.rf._abc_6362_n8403) );
	NAND2X1 NAND2X1_5713 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8403), .Y(dp.rf._abc_6362_n8404) );
	NAND2X1 NAND2X1_5714 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8400), .B(dp.rf._abc_6362_n8404), .Y(dp.rf._abc_6362_n8405) );
	NAND2X1 NAND2X1_5715 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8405), .Y(dp.rf._abc_6362_n8406) );
	NAND2X1 NAND2X1_5716 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8396), .B(dp.rf._abc_6362_n8406), .Y(dp.rf._abc_6362_n8407) );
	NAND2X1 NAND2X1_5717 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n8407), .Y(dp.rf._abc_6362_n8408) );
	NAND2X1 NAND2X1_5718 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n8408), .Y(dp.rf._abc_6362_n8409) );
	NOR2X1 NOR2X1_849 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8386), .B(dp.rf._abc_6362_n8409), .Y(dp.rf._abc_6362_n8410) );
	NAND2X1 NAND2X1_5719 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<30>), .Y(dp.rf._abc_6362_n8411) );
	NAND2X1 NAND2X1_5720 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8412) );
	NAND2X1 NAND2X1_5721 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8411), .B(dp.rf._abc_6362_n8412), .Y(dp.rf._abc_6362_n8413) );
	NAND2X1 NAND2X1_5722 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8413), .Y(dp.rf._abc_6362_n8414) );
	NAND2X1 NAND2X1_5723 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<30>), .Y(dp.rf._abc_6362_n8415) );
	NAND2X1 NAND2X1_5724 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8416) );
	NAND2X1 NAND2X1_5725 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8415), .B(dp.rf._abc_6362_n8416), .Y(dp.rf._abc_6362_n8417) );
	NAND2X1 NAND2X1_5726 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8417), .Y(dp.rf._abc_6362_n8418) );
	AND2X2 AND2X2_329 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8414), .B(dp.rf._abc_6362_n8418), .Y(dp.rf._abc_6362_n8419) );
	NAND2X1 NAND2X1_5727 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8419), .Y(dp.rf._abc_6362_n8420) );
	NAND2X1 NAND2X1_5728 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<30>), .Y(dp.rf._abc_6362_n8421) );
	NAND2X1 NAND2X1_5729 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8422) );
	NAND2X1 NAND2X1_5730 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8421), .B(dp.rf._abc_6362_n8422), .Y(dp.rf._abc_6362_n8423) );
	NAND2X1 NAND2X1_5731 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8423), .Y(dp.rf._abc_6362_n8424) );
	NAND2X1 NAND2X1_5732 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<30>), .Y(dp.rf._abc_6362_n8425) );
	NAND2X1 NAND2X1_5733 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8426) );
	NAND2X1 NAND2X1_5734 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8425), .B(dp.rf._abc_6362_n8426), .Y(dp.rf._abc_6362_n8427) );
	NAND2X1 NAND2X1_5735 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8427), .Y(dp.rf._abc_6362_n8428) );
	AND2X2 AND2X2_330 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8424), .B(dp.rf._abc_6362_n8428), .Y(dp.rf._abc_6362_n8429) );
	NAND2X1 NAND2X1_5736 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8429), .Y(dp.rf._abc_6362_n8430) );
	AND2X2 AND2X2_331 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8430), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n8431) );
	NAND2X1 NAND2X1_5737 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8420), .B(dp.rf._abc_6362_n8431), .Y(dp.rf._abc_6362_n8432) );
	NAND2X1 NAND2X1_5738 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8433) );
	NAND2X1 NAND2X1_5739 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<30>), .Y(dp.rf._abc_6362_n8434) );
	AND2X2 AND2X2_332 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8434), .B(instr[22]), .Y(dp.rf._abc_6362_n8435) );
	NAND2X1 NAND2X1_5740 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8433), .B(dp.rf._abc_6362_n8435), .Y(dp.rf._abc_6362_n8436) );
	NAND2X1 NAND2X1_5741 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8437) );
	NAND2X1 NAND2X1_5742 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<30>), .Y(dp.rf._abc_6362_n8438) );
	AND2X2 AND2X2_333 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8438), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8439) );
	NAND2X1 NAND2X1_5743 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8437), .B(dp.rf._abc_6362_n8439), .Y(dp.rf._abc_6362_n8440) );
	NAND2X1 NAND2X1_5744 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8436), .B(dp.rf._abc_6362_n8440), .Y(dp.rf._abc_6362_n8441) );
	AND2X2 AND2X2_334 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8441), .B(instr[23]), .Y(dp.rf._abc_6362_n8442) );
	NAND2X1 NAND2X1_5745 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8443) );
	NAND2X1 NAND2X1_5746 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<30>), .Y(dp.rf._abc_6362_n8444) );
	AND2X2 AND2X2_335 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8444), .B(instr[22]), .Y(dp.rf._abc_6362_n8445) );
	NAND2X1 NAND2X1_5747 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8443), .B(dp.rf._abc_6362_n8445), .Y(dp.rf._abc_6362_n8446) );
	NAND2X1 NAND2X1_5748 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<30>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8447) );
	NAND2X1 NAND2X1_5749 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<30>), .Y(dp.rf._abc_6362_n8448) );
	AND2X2 AND2X2_336 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8448), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8449) );
	NAND2X1 NAND2X1_5750 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8447), .B(dp.rf._abc_6362_n8449), .Y(dp.rf._abc_6362_n8450) );
	NAND2X1 NAND2X1_5751 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8446), .B(dp.rf._abc_6362_n8450), .Y(dp.rf._abc_6362_n8451) );
	NAND2X1 NAND2X1_5752 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8451), .Y(dp.rf._abc_6362_n8452) );
	NAND2X1 NAND2X1_5753 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n8452), .Y(dp.rf._abc_6362_n8453) );
	NOR2X1 NOR2X1_850 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8442), .B(dp.rf._abc_6362_n8453), .Y(dp.rf._abc_6362_n8454) );
	NOR2X1 NOR2X1_851 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n8454), .Y(dp.rf._abc_6362_n8455) );
	NAND2X1 NAND2X1_5754 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8432), .B(dp.rf._abc_6362_n8455), .Y(dp.rf._abc_6362_n8456) );
	NAND2X1 NAND2X1_5755 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n8456), .Y(dp.rf._abc_6362_n8457) );
	NOR2X1 NOR2X1_852 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8410), .B(dp.rf._abc_6362_n8457), .Y(dp.srca_30_) );
	NAND2X1 NAND2X1_5756 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_11_<31>), .Y(dp.rf._abc_6362_n8459) );
	NAND2X1 NAND2X1_5757 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8459), .Y(dp.rf._abc_6362_n8460) );
	INVX1 INVX1_246 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<31>), .Y(dp.rf._abc_6362_n8461) );
	NOR2X1 NOR2X1_853 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8461), .Y(dp.rf._abc_6362_n8462) );
	NOR2X1 NOR2X1_854 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8460), .B(dp.rf._abc_6362_n8462), .Y(dp.rf._abc_6362_n8463) );
	NAND2X1 NAND2X1_5758 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_9_<31>), .Y(dp.rf._abc_6362_n8464) );
	NAND2X1 NAND2X1_5759 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8464), .Y(dp.rf._abc_6362_n8465) );
	INVX1 INVX1_247 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<31>), .Y(dp.rf._abc_6362_n8466) );
	NOR2X1 NOR2X1_855 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8466), .Y(dp.rf._abc_6362_n8467) );
	NOR2X1 NOR2X1_856 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8465), .B(dp.rf._abc_6362_n8467), .Y(dp.rf._abc_6362_n8468) );
	NOR2X1 NOR2X1_857 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8463), .B(dp.rf._abc_6362_n8468), .Y(dp.rf._abc_6362_n8469) );
	NAND2X1 NAND2X1_5760 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8469), .Y(dp.rf._abc_6362_n8470) );
	NAND2X1 NAND2X1_5761 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_15_<31>), .Y(dp.rf._abc_6362_n8471) );
	NAND2X1 NAND2X1_5762 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8471), .Y(dp.rf._abc_6362_n8472) );
	INVX1 INVX1_248 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<31>), .Y(dp.rf._abc_6362_n8473) );
	NOR2X1 NOR2X1_858 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8473), .Y(dp.rf._abc_6362_n8474) );
	NOR2X1 NOR2X1_859 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8472), .B(dp.rf._abc_6362_n8474), .Y(dp.rf._abc_6362_n8475) );
	NAND2X1 NAND2X1_5763 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_13_<31>), .Y(dp.rf._abc_6362_n8476) );
	NAND2X1 NAND2X1_5764 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8476), .Y(dp.rf._abc_6362_n8477) );
	INVX1 INVX1_249 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<31>), .Y(dp.rf._abc_6362_n8478) );
	NOR2X1 NOR2X1_860 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8478), .Y(dp.rf._abc_6362_n8479) );
	NOR2X1 NOR2X1_861 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8477), .B(dp.rf._abc_6362_n8479), .Y(dp.rf._abc_6362_n8480) );
	NOR2X1 NOR2X1_862 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8475), .B(dp.rf._abc_6362_n8480), .Y(dp.rf._abc_6362_n8481) );
	NAND2X1 NAND2X1_5765 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8481), .Y(dp.rf._abc_6362_n8482) );
	NAND2X1 NAND2X1_5766 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8470), .B(dp.rf._abc_6362_n8482), .Y(dp.rf._abc_6362_n8483) );
	NAND2X1 NAND2X1_5767 ( .gnd(gnd), .vdd(vdd), .A(instr[24]), .B(dp.rf._abc_6362_n8483), .Y(dp.rf._abc_6362_n8484) );
	NAND2X1 NAND2X1_5768 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_7_<31>), .Y(dp.rf._abc_6362_n8485) );
	NAND2X1 NAND2X1_5769 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8485), .Y(dp.rf._abc_6362_n8486) );
	INVX1 INVX1_250 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<31>), .Y(dp.rf._abc_6362_n8487) );
	NOR2X1 NOR2X1_863 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8487), .Y(dp.rf._abc_6362_n8488) );
	NOR2X1 NOR2X1_864 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8486), .B(dp.rf._abc_6362_n8488), .Y(dp.rf._abc_6362_n8489) );
	NAND2X1 NAND2X1_5770 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_5_<31>), .Y(dp.rf._abc_6362_n8490) );
	NAND2X1 NAND2X1_5771 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8490), .Y(dp.rf._abc_6362_n8491) );
	INVX1 INVX1_251 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<31>), .Y(dp.rf._abc_6362_n8492) );
	NOR2X1 NOR2X1_865 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8492), .Y(dp.rf._abc_6362_n8493) );
	NOR2X1 NOR2X1_866 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8491), .B(dp.rf._abc_6362_n8493), .Y(dp.rf._abc_6362_n8494) );
	OR2X2 OR2X2_80 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8489), .B(dp.rf._abc_6362_n8494), .Y(dp.rf._abc_6362_n8495) );
	NAND2X1 NAND2X1_5772 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8495), .Y(dp.rf._abc_6362_n8496) );
	NAND2X1 NAND2X1_5773 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_3_<31>), .Y(dp.rf._abc_6362_n8497) );
	NAND2X1 NAND2X1_5774 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8497), .Y(dp.rf._abc_6362_n8498) );
	INVX1 INVX1_252 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<31>), .Y(dp.rf._abc_6362_n8499) );
	NOR2X1 NOR2X1_867 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8499), .Y(dp.rf._abc_6362_n8500) );
	NOR2X1 NOR2X1_868 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8498), .B(dp.rf._abc_6362_n8500), .Y(dp.rf._abc_6362_n8501) );
	NAND2X1 NAND2X1_5775 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_1_<31>), .Y(dp.rf._abc_6362_n8502) );
	NAND2X1 NAND2X1_5776 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8502), .Y(dp.rf._abc_6362_n8503) );
	INVX1 INVX1_253 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<31>), .Y(dp.rf._abc_6362_n8504) );
	NOR2X1 NOR2X1_869 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf._abc_6362_n8504), .Y(dp.rf._abc_6362_n8505) );
	NOR2X1 NOR2X1_870 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8503), .B(dp.rf._abc_6362_n8505), .Y(dp.rf._abc_6362_n8506) );
	OR2X2 OR2X2_81 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8501), .B(dp.rf._abc_6362_n8506), .Y(dp.rf._abc_6362_n8507) );
	NAND2X1 NAND2X1_5777 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8507), .Y(dp.rf._abc_6362_n8508) );
	AND2X2 AND2X2_337 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8508), .B(dp.rf._abc_6362_n5397), .Y(dp.rf._abc_6362_n8509) );
	NAND2X1 NAND2X1_5778 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8496), .B(dp.rf._abc_6362_n8509), .Y(dp.rf._abc_6362_n8510) );
	NAND2X1 NAND2X1_5779 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8484), .B(dp.rf._abc_6362_n8510), .Y(dp.rf._abc_6362_n8511) );
	NOR2X1 NOR2X1_871 ( .gnd(gnd), .vdd(vdd), .A(instr[25]), .B(dp.rf._abc_6362_n8511), .Y(dp.rf._abc_6362_n8512) );
	NAND2X1 NAND2X1_5780 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_25_<31>), .Y(dp.rf._abc_6362_n8513) );
	NAND2X1 NAND2X1_5781 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<31>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8514) );
	NAND2X1 NAND2X1_5782 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8513), .B(dp.rf._abc_6362_n8514), .Y(dp.rf._abc_6362_n8515) );
	NAND2X1 NAND2X1_5783 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8515), .Y(dp.rf._abc_6362_n8516) );
	NAND2X1 NAND2X1_5784 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_27_<31>), .Y(dp.rf._abc_6362_n8517) );
	NAND2X1 NAND2X1_5785 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<31>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8518) );
	NAND2X1 NAND2X1_5786 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8517), .B(dp.rf._abc_6362_n8518), .Y(dp.rf._abc_6362_n8519) );
	NAND2X1 NAND2X1_5787 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8519), .Y(dp.rf._abc_6362_n8520) );
	AND2X2 AND2X2_338 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8516), .B(dp.rf._abc_6362_n8520), .Y(dp.rf._abc_6362_n8521) );
	NAND2X1 NAND2X1_5788 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8521), .Y(dp.rf._abc_6362_n8522) );
	NAND2X1 NAND2X1_5789 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_29_<31>), .Y(dp.rf._abc_6362_n8523) );
	NAND2X1 NAND2X1_5790 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<31>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8524) );
	NAND2X1 NAND2X1_5791 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8523), .B(dp.rf._abc_6362_n8524), .Y(dp.rf._abc_6362_n8525) );
	NAND2X1 NAND2X1_5792 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5340), .B(dp.rf._abc_6362_n8525), .Y(dp.rf._abc_6362_n8526) );
	NAND2X1 NAND2X1_5793 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_31_<31>), .Y(dp.rf._abc_6362_n8527) );
	NAND2X1 NAND2X1_5794 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<31>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8528) );
	NAND2X1 NAND2X1_5795 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8527), .B(dp.rf._abc_6362_n8528), .Y(dp.rf._abc_6362_n8529) );
	NAND2X1 NAND2X1_5796 ( .gnd(gnd), .vdd(vdd), .A(instr[22]), .B(dp.rf._abc_6362_n8529), .Y(dp.rf._abc_6362_n8530) );
	AND2X2 AND2X2_339 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8526), .B(dp.rf._abc_6362_n8530), .Y(dp.rf._abc_6362_n8531) );
	NAND2X1 NAND2X1_5797 ( .gnd(gnd), .vdd(vdd), .A(instr[23]), .B(dp.rf._abc_6362_n8531), .Y(dp.rf._abc_6362_n8532) );
	AND2X2 AND2X2_340 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8532), .B(instr[24]), .Y(dp.rf._abc_6362_n8533) );
	NAND2X1 NAND2X1_5798 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8522), .B(dp.rf._abc_6362_n8533), .Y(dp.rf._abc_6362_n8534) );
	NAND2X1 NAND2X1_5799 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<31>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8535) );
	NAND2X1 NAND2X1_5800 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_23_<31>), .Y(dp.rf._abc_6362_n8536) );
	AND2X2 AND2X2_341 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8536), .B(instr[22]), .Y(dp.rf._abc_6362_n8537) );
	NAND2X1 NAND2X1_5801 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8535), .B(dp.rf._abc_6362_n8537), .Y(dp.rf._abc_6362_n8538) );
	NAND2X1 NAND2X1_5802 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<31>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8539) );
	NAND2X1 NAND2X1_5803 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_21_<31>), .Y(dp.rf._abc_6362_n8540) );
	AND2X2 AND2X2_342 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8540), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8541) );
	NAND2X1 NAND2X1_5804 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8539), .B(dp.rf._abc_6362_n8541), .Y(dp.rf._abc_6362_n8542) );
	NAND2X1 NAND2X1_5805 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8538), .B(dp.rf._abc_6362_n8542), .Y(dp.rf._abc_6362_n8543) );
	AND2X2 AND2X2_343 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8543), .B(instr[23]), .Y(dp.rf._abc_6362_n8544) );
	NAND2X1 NAND2X1_5806 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<31>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8545) );
	NAND2X1 NAND2X1_5807 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_19_<31>), .Y(dp.rf._abc_6362_n8546) );
	AND2X2 AND2X2_344 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8546), .B(instr[22]), .Y(dp.rf._abc_6362_n8547) );
	NAND2X1 NAND2X1_5808 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8545), .B(dp.rf._abc_6362_n8547), .Y(dp.rf._abc_6362_n8548) );
	NAND2X1 NAND2X1_5809 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<31>), .B(dp.rf._abc_6362_n5338), .Y(dp.rf._abc_6362_n8549) );
	NAND2X1 NAND2X1_5810 ( .gnd(gnd), .vdd(vdd), .A(instr[21]), .B(dp.rf.rf_17_<31>), .Y(dp.rf._abc_6362_n8550) );
	AND2X2 AND2X2_345 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8550), .B(dp.rf._abc_6362_n5340), .Y(dp.rf._abc_6362_n8551) );
	NAND2X1 NAND2X1_5811 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8549), .B(dp.rf._abc_6362_n8551), .Y(dp.rf._abc_6362_n8552) );
	NAND2X1 NAND2X1_5812 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8548), .B(dp.rf._abc_6362_n8552), .Y(dp.rf._abc_6362_n8553) );
	NAND2X1 NAND2X1_5813 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5352), .B(dp.rf._abc_6362_n8553), .Y(dp.rf._abc_6362_n8554) );
	NAND2X1 NAND2X1_5814 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5397), .B(dp.rf._abc_6362_n8554), .Y(dp.rf._abc_6362_n8555) );
	NOR2X1 NOR2X1_872 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8544), .B(dp.rf._abc_6362_n8555), .Y(dp.rf._abc_6362_n8556) );
	NOR2X1 NOR2X1_873 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5367), .B(dp.rf._abc_6362_n8556), .Y(dp.rf._abc_6362_n8557) );
	NAND2X1 NAND2X1_5815 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8534), .B(dp.rf._abc_6362_n8557), .Y(dp.rf._abc_6362_n8558) );
	NAND2X1 NAND2X1_5816 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n5400), .B(dp.rf._abc_6362_n8558), .Y(dp.rf._abc_6362_n8559) );
	NOR2X1 NOR2X1_874 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8512), .B(dp.rf._abc_6362_n8559), .Y(dp.srca_31_) );
	INVX8 INVX8_42 ( .gnd(gnd), .vdd(vdd), .A(instr[20]), .Y(dp.rf._abc_6362_n8561) );
	INVX8 INVX8_43 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .Y(dp.rf._abc_6362_n8562) );
	NAND2X1 NAND2X1_5817 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<0>), .Y(dp.rf._abc_6362_n8563) );
	NAND2X1 NAND2X1_5818 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8563), .Y(dp.rf._abc_6362_n8564) );
	NOR2X1 NOR2X1_875 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5382), .Y(dp.rf._abc_6362_n8565) );
	NOR2X1 NOR2X1_876 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8564), .B(dp.rf._abc_6362_n8565), .Y(dp.rf._abc_6362_n8566) );
	INVX8 INVX8_44 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .Y(dp.rf._abc_6362_n8567) );
	NAND2X1 NAND2X1_5819 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<0>), .Y(dp.rf._abc_6362_n8568) );
	NAND2X1 NAND2X1_5820 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8568), .Y(dp.rf._abc_6362_n8569) );
	NOR2X1 NOR2X1_877 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5387), .Y(dp.rf._abc_6362_n8570) );
	NOR2X1 NOR2X1_878 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8569), .B(dp.rf._abc_6362_n8570), .Y(dp.rf._abc_6362_n8571) );
	NOR2X1 NOR2X1_879 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8566), .B(dp.rf._abc_6362_n8571), .Y(dp.rf._abc_6362_n8572) );
	NAND2X1 NAND2X1_5821 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8572), .Y(dp.rf._abc_6362_n8573) );
	NAND2X1 NAND2X1_5822 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<0>), .Y(dp.rf._abc_6362_n8574) );
	NAND2X1 NAND2X1_5823 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8574), .Y(dp.rf._abc_6362_n8575) );
	NOR2X1 NOR2X1_880 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5370), .Y(dp.rf._abc_6362_n8576) );
	NOR2X1 NOR2X1_881 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8575), .B(dp.rf._abc_6362_n8576), .Y(dp.rf._abc_6362_n8577) );
	NAND2X1 NAND2X1_5824 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<0>), .Y(dp.rf._abc_6362_n8578) );
	NAND2X1 NAND2X1_5825 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8578), .Y(dp.rf._abc_6362_n8579) );
	NOR2X1 NOR2X1_882 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5375), .Y(dp.rf._abc_6362_n8580) );
	NOR2X1 NOR2X1_883 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8579), .B(dp.rf._abc_6362_n8580), .Y(dp.rf._abc_6362_n8581) );
	NOR2X1 NOR2X1_884 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8577), .B(dp.rf._abc_6362_n8581), .Y(dp.rf._abc_6362_n8582) );
	NAND2X1 NAND2X1_5826 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8582), .Y(dp.rf._abc_6362_n8583) );
	NAND2X1 NAND2X1_5827 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8573), .B(dp.rf._abc_6362_n8583), .Y(dp.rf._abc_6362_n8584) );
	NAND2X1 NAND2X1_5828 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n8584), .Y(dp.rf._abc_6362_n8585) );
	NAND2X1 NAND2X1_5829 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n8585), .Y(dp.rf._abc_6362_n8586) );
	INVX8 INVX8_45 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .Y(dp.rf._abc_6362_n8587) );
	NAND2X1 NAND2X1_5830 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<0>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8588) );
	NOR2X1 NOR2X1_885 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5354), .Y(dp.rf._abc_6362_n8589) );
	NOR2X1 NOR2X1_886 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8589), .Y(dp.rf._abc_6362_n8590) );
	NAND2X1 NAND2X1_5831 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8588), .B(dp.rf._abc_6362_n8590), .Y(dp.rf._abc_6362_n8591) );
	NAND2X1 NAND2X1_5832 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<0>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8592) );
	NOR2X1 NOR2X1_887 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5359), .Y(dp.rf._abc_6362_n8593) );
	NOR2X1 NOR2X1_888 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8593), .Y(dp.rf._abc_6362_n8594) );
	NAND2X1 NAND2X1_5833 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8592), .B(dp.rf._abc_6362_n8594), .Y(dp.rf._abc_6362_n8595) );
	NAND2X1 NAND2X1_5834 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8591), .B(dp.rf._abc_6362_n8595), .Y(dp.rf._abc_6362_n8596) );
	NOR2X1 NOR2X1_889 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8596), .Y(dp.rf._abc_6362_n8597) );
	NAND2X1 NAND2X1_5835 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<0>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8598) );
	NOR2X1 NOR2X1_890 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5341), .Y(dp.rf._abc_6362_n8599) );
	NOR2X1 NOR2X1_891 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8599), .Y(dp.rf._abc_6362_n8600) );
	NAND2X1 NAND2X1_5836 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8598), .B(dp.rf._abc_6362_n8600), .Y(dp.rf._abc_6362_n8601) );
	NAND2X1 NAND2X1_5837 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<0>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8602) );
	NOR2X1 NOR2X1_892 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5346), .Y(dp.rf._abc_6362_n8603) );
	NOR2X1 NOR2X1_893 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8603), .Y(dp.rf._abc_6362_n8604) );
	NAND2X1 NAND2X1_5838 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8602), .B(dp.rf._abc_6362_n8604), .Y(dp.rf._abc_6362_n8605) );
	NAND2X1 NAND2X1_5839 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8601), .B(dp.rf._abc_6362_n8605), .Y(dp.rf._abc_6362_n8606) );
	NOR2X1 NOR2X1_894 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8606), .Y(dp.rf._abc_6362_n8607) );
	NOR2X1 NOR2X1_895 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8597), .B(dp.rf._abc_6362_n8607), .Y(dp.rf._abc_6362_n8608) );
	NOR2X1 NOR2X1_896 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n8608), .Y(dp.rf._abc_6362_n8609) );
	NOR2X1 NOR2X1_897 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8586), .B(dp.rf._abc_6362_n8609), .Y(dp.rf._abc_6362_n8610) );
	NOR2X1 NOR2X1_898 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(instr[17]), .Y(dp.rf._abc_6362_n8611) );
	INVX8 INVX8_46 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .Y(dp.rf._abc_6362_n8612) );
	NAND2X1 NAND2X1_5840 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n8613) );
	NOR2X1 NOR2X1_899 ( .gnd(gnd), .vdd(vdd), .A(instr[20]), .B(dp.rf._abc_6362_n8613), .Y(dp.rf._abc_6362_n8614) );
	NAND2X1 NAND2X1_5841 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8611), .B(dp.rf._abc_6362_n8614), .Y(dp.rf._abc_6362_n8615) );
	NAND2X1 NAND2X1_5842 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<0>), .Y(dp.rf._abc_6362_n8616) );
	NAND2X1 NAND2X1_5843 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8616), .Y(dp.rf._abc_6362_n8617) );
	NOR2X1 NOR2X1_900 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5403), .Y(dp.rf._abc_6362_n8618) );
	NOR2X1 NOR2X1_901 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8617), .B(dp.rf._abc_6362_n8618), .Y(dp.rf._abc_6362_n8619) );
	NAND2X1 NAND2X1_5844 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<0>), .Y(dp.rf._abc_6362_n8620) );
	NAND2X1 NAND2X1_5845 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8620), .Y(dp.rf._abc_6362_n8621) );
	NOR2X1 NOR2X1_902 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5408), .Y(dp.rf._abc_6362_n8622) );
	NOR2X1 NOR2X1_903 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8621), .B(dp.rf._abc_6362_n8622), .Y(dp.rf._abc_6362_n8623) );
	OR2X2 OR2X2_82 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8619), .B(dp.rf._abc_6362_n8623), .Y(dp.rf._abc_6362_n8624) );
	NAND2X1 NAND2X1_5846 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8624), .Y(dp.rf._abc_6362_n8625) );
	NAND2X1 NAND2X1_5847 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<0>), .Y(dp.rf._abc_6362_n8626) );
	NAND2X1 NAND2X1_5848 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8626), .Y(dp.rf._abc_6362_n8627) );
	NOR2X1 NOR2X1_904 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5415), .Y(dp.rf._abc_6362_n8628) );
	NOR2X1 NOR2X1_905 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8627), .B(dp.rf._abc_6362_n8628), .Y(dp.rf._abc_6362_n8629) );
	NAND2X1 NAND2X1_5849 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<0>), .Y(dp.rf._abc_6362_n8630) );
	NAND2X1 NAND2X1_5850 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8630), .Y(dp.rf._abc_6362_n8631) );
	NOR2X1 NOR2X1_906 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5420), .Y(dp.rf._abc_6362_n8632) );
	NOR2X1 NOR2X1_907 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8631), .B(dp.rf._abc_6362_n8632), .Y(dp.rf._abc_6362_n8633) );
	OR2X2 OR2X2_83 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8629), .B(dp.rf._abc_6362_n8633), .Y(dp.rf._abc_6362_n8634) );
	NAND2X1 NAND2X1_5851 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8634), .Y(dp.rf._abc_6362_n8635) );
	AND2X2 AND2X2_346 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8635), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n8636) );
	NAND2X1 NAND2X1_5852 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8625), .B(dp.rf._abc_6362_n8636), .Y(dp.rf._abc_6362_n8637) );
	NAND2X1 NAND2X1_5853 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<0>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8638) );
	NAND2X1 NAND2X1_5854 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<0>), .Y(dp.rf._abc_6362_n8639) );
	AND2X2 AND2X2_347 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8639), .B(instr[17]), .Y(dp.rf._abc_6362_n8640) );
	NAND2X1 NAND2X1_5855 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8638), .B(dp.rf._abc_6362_n8640), .Y(dp.rf._abc_6362_n8641) );
	NAND2X1 NAND2X1_5856 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<0>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8642) );
	NAND2X1 NAND2X1_5857 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<0>), .Y(dp.rf._abc_6362_n8643) );
	AND2X2 AND2X2_348 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8643), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n8644) );
	NAND2X1 NAND2X1_5858 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8642), .B(dp.rf._abc_6362_n8644), .Y(dp.rf._abc_6362_n8645) );
	NAND2X1 NAND2X1_5859 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8641), .B(dp.rf._abc_6362_n8645), .Y(dp.rf._abc_6362_n8646) );
	AND2X2 AND2X2_349 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8646), .B(instr[18]), .Y(dp.rf._abc_6362_n8647) );
	NAND2X1 NAND2X1_5860 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<0>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8648) );
	NAND2X1 NAND2X1_5861 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<0>), .Y(dp.rf._abc_6362_n8649) );
	AND2X2 AND2X2_350 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8649), .B(instr[17]), .Y(dp.rf._abc_6362_n8650) );
	NAND2X1 NAND2X1_5862 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8648), .B(dp.rf._abc_6362_n8650), .Y(dp.rf._abc_6362_n8651) );
	NAND2X1 NAND2X1_5863 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<0>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8652) );
	NAND2X1 NAND2X1_5864 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<0>), .Y(dp.rf._abc_6362_n8653) );
	AND2X2 AND2X2_351 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8653), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n8654) );
	NAND2X1 NAND2X1_5865 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8652), .B(dp.rf._abc_6362_n8654), .Y(dp.rf._abc_6362_n8655) );
	NAND2X1 NAND2X1_5866 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8651), .B(dp.rf._abc_6362_n8655), .Y(dp.rf._abc_6362_n8656) );
	NAND2X1 NAND2X1_5867 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8656), .Y(dp.rf._abc_6362_n8657) );
	NAND2X1 NAND2X1_5868 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n8657), .Y(dp.rf._abc_6362_n8658) );
	NOR2X1 NOR2X1_908 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8647), .B(dp.rf._abc_6362_n8658), .Y(dp.rf._abc_6362_n8659) );
	NOR2X1 NOR2X1_909 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n8659), .Y(dp.rf._abc_6362_n8660) );
	NAND2X1 NAND2X1_5869 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8637), .B(dp.rf._abc_6362_n8660), .Y(dp.rf._abc_6362_n8661) );
	NAND2X1 NAND2X1_5870 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n8661), .Y(dp.rf._abc_6362_n8662) );
	NOR2X1 NOR2X1_910 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8610), .B(dp.rf._abc_6362_n8662), .Y(writedata_0__RAW) );
	NAND2X1 NAND2X1_5871 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8664) );
	NOR2X1 NOR2X1_911 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5481), .Y(dp.rf._abc_6362_n8665) );
	NOR2X1 NOR2X1_912 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8665), .Y(dp.rf._abc_6362_n8666) );
	NAND2X1 NAND2X1_5872 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8664), .B(dp.rf._abc_6362_n8666), .Y(dp.rf._abc_6362_n8667) );
	NAND2X1 NAND2X1_5873 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8668) );
	NOR2X1 NOR2X1_913 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5486), .Y(dp.rf._abc_6362_n8669) );
	NOR2X1 NOR2X1_914 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8669), .Y(dp.rf._abc_6362_n8670) );
	NAND2X1 NAND2X1_5874 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8668), .B(dp.rf._abc_6362_n8670), .Y(dp.rf._abc_6362_n8671) );
	NAND2X1 NAND2X1_5875 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8667), .B(dp.rf._abc_6362_n8671), .Y(dp.rf._abc_6362_n8672) );
	NOR2X1 NOR2X1_915 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8672), .Y(dp.rf._abc_6362_n8673) );
	NAND2X1 NAND2X1_5876 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8674) );
	NOR2X1 NOR2X1_916 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5493), .Y(dp.rf._abc_6362_n8675) );
	NOR2X1 NOR2X1_917 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8675), .Y(dp.rf._abc_6362_n8676) );
	NAND2X1 NAND2X1_5877 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8674), .B(dp.rf._abc_6362_n8676), .Y(dp.rf._abc_6362_n8677) );
	NAND2X1 NAND2X1_5878 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8678) );
	NOR2X1 NOR2X1_918 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5498), .Y(dp.rf._abc_6362_n8679) );
	NOR2X1 NOR2X1_919 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8679), .Y(dp.rf._abc_6362_n8680) );
	NAND2X1 NAND2X1_5879 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8678), .B(dp.rf._abc_6362_n8680), .Y(dp.rf._abc_6362_n8681) );
	NAND2X1 NAND2X1_5880 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8677), .B(dp.rf._abc_6362_n8681), .Y(dp.rf._abc_6362_n8682) );
	NOR2X1 NOR2X1_920 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8682), .Y(dp.rf._abc_6362_n8683) );
	NOR2X1 NOR2X1_921 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8673), .B(dp.rf._abc_6362_n8683), .Y(dp.rf._abc_6362_n8684) );
	NOR2X1 NOR2X1_922 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n8684), .Y(dp.rf._abc_6362_n8685) );
	NAND2X1 NAND2X1_5881 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<1>), .Y(dp.rf._abc_6362_n8686) );
	NAND2X1 NAND2X1_5882 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8686), .Y(dp.rf._abc_6362_n8687) );
	NOR2X1 NOR2X1_923 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5467), .Y(dp.rf._abc_6362_n8688) );
	NOR2X1 NOR2X1_924 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8687), .B(dp.rf._abc_6362_n8688), .Y(dp.rf._abc_6362_n8689) );
	NAND2X1 NAND2X1_5883 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<1>), .Y(dp.rf._abc_6362_n8690) );
	NAND2X1 NAND2X1_5884 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8690), .Y(dp.rf._abc_6362_n8691) );
	NOR2X1 NOR2X1_925 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5472), .Y(dp.rf._abc_6362_n8692) );
	NOR2X1 NOR2X1_926 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8691), .B(dp.rf._abc_6362_n8692), .Y(dp.rf._abc_6362_n8693) );
	OR2X2 OR2X2_84 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8689), .B(dp.rf._abc_6362_n8693), .Y(dp.rf._abc_6362_n8694) );
	NAND2X1 NAND2X1_5885 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8694), .Y(dp.rf._abc_6362_n8695) );
	NAND2X1 NAND2X1_5886 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<1>), .Y(dp.rf._abc_6362_n8696) );
	NAND2X1 NAND2X1_5887 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8696), .Y(dp.rf._abc_6362_n8697) );
	NOR2X1 NOR2X1_927 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5455), .Y(dp.rf._abc_6362_n8698) );
	NOR2X1 NOR2X1_928 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8697), .B(dp.rf._abc_6362_n8698), .Y(dp.rf._abc_6362_n8699) );
	NAND2X1 NAND2X1_5888 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<1>), .Y(dp.rf._abc_6362_n8700) );
	NAND2X1 NAND2X1_5889 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8700), .Y(dp.rf._abc_6362_n8701) );
	NOR2X1 NOR2X1_929 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5460), .Y(dp.rf._abc_6362_n8702) );
	NOR2X1 NOR2X1_930 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8701), .B(dp.rf._abc_6362_n8702), .Y(dp.rf._abc_6362_n8703) );
	OR2X2 OR2X2_85 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8699), .B(dp.rf._abc_6362_n8703), .Y(dp.rf._abc_6362_n8704) );
	NAND2X1 NAND2X1_5890 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8704), .Y(dp.rf._abc_6362_n8705) );
	AND2X2 AND2X2_352 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8705), .B(instr[19]), .Y(dp.rf._abc_6362_n8706) );
	NAND2X1 NAND2X1_5891 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8695), .B(dp.rf._abc_6362_n8706), .Y(dp.rf._abc_6362_n8707) );
	NAND2X1 NAND2X1_5892 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n8707), .Y(dp.rf._abc_6362_n8708) );
	NOR2X1 NOR2X1_931 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8685), .B(dp.rf._abc_6362_n8708), .Y(dp.rf._abc_6362_n8709) );
	NAND2X1 NAND2X1_5893 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<1>), .Y(dp.rf._abc_6362_n8710) );
	NAND2X1 NAND2X1_5894 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8711) );
	NAND2X1 NAND2X1_5895 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8710), .B(dp.rf._abc_6362_n8711), .Y(dp.rf._abc_6362_n8712) );
	NAND2X1 NAND2X1_5896 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8712), .Y(dp.rf._abc_6362_n8713) );
	NAND2X1 NAND2X1_5897 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<1>), .Y(dp.rf._abc_6362_n8714) );
	NAND2X1 NAND2X1_5898 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8715) );
	NAND2X1 NAND2X1_5899 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8714), .B(dp.rf._abc_6362_n8715), .Y(dp.rf._abc_6362_n8716) );
	NAND2X1 NAND2X1_5900 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8716), .Y(dp.rf._abc_6362_n8717) );
	AND2X2 AND2X2_353 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8713), .B(dp.rf._abc_6362_n8717), .Y(dp.rf._abc_6362_n8718) );
	NAND2X1 NAND2X1_5901 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8718), .Y(dp.rf._abc_6362_n8719) );
	NAND2X1 NAND2X1_5902 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<1>), .Y(dp.rf._abc_6362_n8720) );
	NAND2X1 NAND2X1_5903 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8721) );
	NAND2X1 NAND2X1_5904 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8720), .B(dp.rf._abc_6362_n8721), .Y(dp.rf._abc_6362_n8722) );
	NAND2X1 NAND2X1_5905 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8722), .Y(dp.rf._abc_6362_n8723) );
	NAND2X1 NAND2X1_5906 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<1>), .Y(dp.rf._abc_6362_n8724) );
	NAND2X1 NAND2X1_5907 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8725) );
	NAND2X1 NAND2X1_5908 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8724), .B(dp.rf._abc_6362_n8725), .Y(dp.rf._abc_6362_n8726) );
	NAND2X1 NAND2X1_5909 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8726), .Y(dp.rf._abc_6362_n8727) );
	AND2X2 AND2X2_354 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8723), .B(dp.rf._abc_6362_n8727), .Y(dp.rf._abc_6362_n8728) );
	NAND2X1 NAND2X1_5910 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8728), .Y(dp.rf._abc_6362_n8729) );
	AND2X2 AND2X2_355 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8729), .B(instr[19]), .Y(dp.rf._abc_6362_n8730) );
	NAND2X1 NAND2X1_5911 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8719), .B(dp.rf._abc_6362_n8730), .Y(dp.rf._abc_6362_n8731) );
	NAND2X1 NAND2X1_5912 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8732) );
	NAND2X1 NAND2X1_5913 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<1>), .Y(dp.rf._abc_6362_n8733) );
	AND2X2 AND2X2_356 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8733), .B(instr[17]), .Y(dp.rf._abc_6362_n8734) );
	NAND2X1 NAND2X1_5914 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8732), .B(dp.rf._abc_6362_n8734), .Y(dp.rf._abc_6362_n8735) );
	NAND2X1 NAND2X1_5915 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8736) );
	NAND2X1 NAND2X1_5916 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<1>), .Y(dp.rf._abc_6362_n8737) );
	AND2X2 AND2X2_357 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8737), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n8738) );
	NAND2X1 NAND2X1_5917 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8736), .B(dp.rf._abc_6362_n8738), .Y(dp.rf._abc_6362_n8739) );
	NAND2X1 NAND2X1_5918 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8735), .B(dp.rf._abc_6362_n8739), .Y(dp.rf._abc_6362_n8740) );
	AND2X2 AND2X2_358 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8740), .B(instr[18]), .Y(dp.rf._abc_6362_n8741) );
	NAND2X1 NAND2X1_5919 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8742) );
	NAND2X1 NAND2X1_5920 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<1>), .Y(dp.rf._abc_6362_n8743) );
	AND2X2 AND2X2_359 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8743), .B(instr[17]), .Y(dp.rf._abc_6362_n8744) );
	NAND2X1 NAND2X1_5921 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8742), .B(dp.rf._abc_6362_n8744), .Y(dp.rf._abc_6362_n8745) );
	NAND2X1 NAND2X1_5922 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<1>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8746) );
	NAND2X1 NAND2X1_5923 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<1>), .Y(dp.rf._abc_6362_n8747) );
	AND2X2 AND2X2_360 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8747), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n8748) );
	NAND2X1 NAND2X1_5924 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8746), .B(dp.rf._abc_6362_n8748), .Y(dp.rf._abc_6362_n8749) );
	NAND2X1 NAND2X1_5925 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8745), .B(dp.rf._abc_6362_n8749), .Y(dp.rf._abc_6362_n8750) );
	NAND2X1 NAND2X1_5926 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8750), .Y(dp.rf._abc_6362_n8751) );
	NAND2X1 NAND2X1_5927 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n8751), .Y(dp.rf._abc_6362_n8752) );
	NOR2X1 NOR2X1_932 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8741), .B(dp.rf._abc_6362_n8752), .Y(dp.rf._abc_6362_n8753) );
	NOR2X1 NOR2X1_933 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n8753), .Y(dp.rf._abc_6362_n8754) );
	NAND2X1 NAND2X1_5928 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8731), .B(dp.rf._abc_6362_n8754), .Y(dp.rf._abc_6362_n8755) );
	NAND2X1 NAND2X1_5929 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n8755), .Y(dp.rf._abc_6362_n8756) );
	NOR2X1 NOR2X1_934 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8709), .B(dp.rf._abc_6362_n8756), .Y(writedata_1__RAW) );
	NAND2X1 NAND2X1_5930 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<2>), .Y(dp.rf._abc_6362_n8758) );
	NAND2X1 NAND2X1_5931 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8758), .Y(dp.rf._abc_6362_n8759) );
	NOR2X1 NOR2X1_935 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5557), .Y(dp.rf._abc_6362_n8760) );
	NOR2X1 NOR2X1_936 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8759), .B(dp.rf._abc_6362_n8760), .Y(dp.rf._abc_6362_n8761) );
	NAND2X1 NAND2X1_5932 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<2>), .Y(dp.rf._abc_6362_n8762) );
	NAND2X1 NAND2X1_5933 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8762), .Y(dp.rf._abc_6362_n8763) );
	NOR2X1 NOR2X1_937 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5562), .Y(dp.rf._abc_6362_n8764) );
	NOR2X1 NOR2X1_938 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8763), .B(dp.rf._abc_6362_n8764), .Y(dp.rf._abc_6362_n8765) );
	NOR2X1 NOR2X1_939 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8761), .B(dp.rf._abc_6362_n8765), .Y(dp.rf._abc_6362_n8766) );
	NAND2X1 NAND2X1_5934 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8766), .Y(dp.rf._abc_6362_n8767) );
	NAND2X1 NAND2X1_5935 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<2>), .Y(dp.rf._abc_6362_n8768) );
	NAND2X1 NAND2X1_5936 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8768), .Y(dp.rf._abc_6362_n8769) );
	NOR2X1 NOR2X1_940 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5569), .Y(dp.rf._abc_6362_n8770) );
	NOR2X1 NOR2X1_941 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8769), .B(dp.rf._abc_6362_n8770), .Y(dp.rf._abc_6362_n8771) );
	NAND2X1 NAND2X1_5937 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<2>), .Y(dp.rf._abc_6362_n8772) );
	NAND2X1 NAND2X1_5938 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8772), .Y(dp.rf._abc_6362_n8773) );
	NOR2X1 NOR2X1_942 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5574), .Y(dp.rf._abc_6362_n8774) );
	NOR2X1 NOR2X1_943 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8773), .B(dp.rf._abc_6362_n8774), .Y(dp.rf._abc_6362_n8775) );
	NOR2X1 NOR2X1_944 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8771), .B(dp.rf._abc_6362_n8775), .Y(dp.rf._abc_6362_n8776) );
	NAND2X1 NAND2X1_5939 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8776), .Y(dp.rf._abc_6362_n8777) );
	NAND2X1 NAND2X1_5940 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8767), .B(dp.rf._abc_6362_n8777), .Y(dp.rf._abc_6362_n8778) );
	NAND2X1 NAND2X1_5941 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n8778), .Y(dp.rf._abc_6362_n8779) );
	NAND2X1 NAND2X1_5942 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n8779), .Y(dp.rf._abc_6362_n8780) );
	NAND2X1 NAND2X1_5943 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8781) );
	NOR2X1 NOR2X1_945 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5583), .Y(dp.rf._abc_6362_n8782) );
	NOR2X1 NOR2X1_946 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8782), .Y(dp.rf._abc_6362_n8783) );
	NAND2X1 NAND2X1_5944 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8781), .B(dp.rf._abc_6362_n8783), .Y(dp.rf._abc_6362_n8784) );
	NAND2X1 NAND2X1_5945 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8785) );
	NOR2X1 NOR2X1_947 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5588), .Y(dp.rf._abc_6362_n8786) );
	NOR2X1 NOR2X1_948 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8786), .Y(dp.rf._abc_6362_n8787) );
	NAND2X1 NAND2X1_5946 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8785), .B(dp.rf._abc_6362_n8787), .Y(dp.rf._abc_6362_n8788) );
	NAND2X1 NAND2X1_5947 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8784), .B(dp.rf._abc_6362_n8788), .Y(dp.rf._abc_6362_n8789) );
	NOR2X1 NOR2X1_949 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8789), .Y(dp.rf._abc_6362_n8790) );
	NAND2X1 NAND2X1_5948 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8791) );
	NOR2X1 NOR2X1_950 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5595), .Y(dp.rf._abc_6362_n8792) );
	NOR2X1 NOR2X1_951 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8792), .Y(dp.rf._abc_6362_n8793) );
	NAND2X1 NAND2X1_5949 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8791), .B(dp.rf._abc_6362_n8793), .Y(dp.rf._abc_6362_n8794) );
	NAND2X1 NAND2X1_5950 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8795) );
	NOR2X1 NOR2X1_952 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5600), .Y(dp.rf._abc_6362_n8796) );
	NOR2X1 NOR2X1_953 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8796), .Y(dp.rf._abc_6362_n8797) );
	NAND2X1 NAND2X1_5951 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8795), .B(dp.rf._abc_6362_n8797), .Y(dp.rf._abc_6362_n8798) );
	NAND2X1 NAND2X1_5952 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8794), .B(dp.rf._abc_6362_n8798), .Y(dp.rf._abc_6362_n8799) );
	NOR2X1 NOR2X1_954 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8799), .Y(dp.rf._abc_6362_n8800) );
	NOR2X1 NOR2X1_955 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8790), .B(dp.rf._abc_6362_n8800), .Y(dp.rf._abc_6362_n8801) );
	NOR2X1 NOR2X1_956 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n8801), .Y(dp.rf._abc_6362_n8802) );
	NOR2X1 NOR2X1_957 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8780), .B(dp.rf._abc_6362_n8802), .Y(dp.rf._abc_6362_n8803) );
	NAND2X1 NAND2X1_5953 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<2>), .Y(dp.rf._abc_6362_n8804) );
	NAND2X1 NAND2X1_5954 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8805) );
	NAND2X1 NAND2X1_5955 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8804), .B(dp.rf._abc_6362_n8805), .Y(dp.rf._abc_6362_n8806) );
	NAND2X1 NAND2X1_5956 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8806), .Y(dp.rf._abc_6362_n8807) );
	NAND2X1 NAND2X1_5957 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<2>), .Y(dp.rf._abc_6362_n8808) );
	NAND2X1 NAND2X1_5958 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8809) );
	NAND2X1 NAND2X1_5959 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8808), .B(dp.rf._abc_6362_n8809), .Y(dp.rf._abc_6362_n8810) );
	NAND2X1 NAND2X1_5960 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8810), .Y(dp.rf._abc_6362_n8811) );
	AND2X2 AND2X2_361 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8807), .B(dp.rf._abc_6362_n8811), .Y(dp.rf._abc_6362_n8812) );
	NAND2X1 NAND2X1_5961 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8812), .Y(dp.rf._abc_6362_n8813) );
	NAND2X1 NAND2X1_5962 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<2>), .Y(dp.rf._abc_6362_n8814) );
	NAND2X1 NAND2X1_5963 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8815) );
	NAND2X1 NAND2X1_5964 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8814), .B(dp.rf._abc_6362_n8815), .Y(dp.rf._abc_6362_n8816) );
	NAND2X1 NAND2X1_5965 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8816), .Y(dp.rf._abc_6362_n8817) );
	NAND2X1 NAND2X1_5966 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<2>), .Y(dp.rf._abc_6362_n8818) );
	NAND2X1 NAND2X1_5967 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8819) );
	NAND2X1 NAND2X1_5968 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8818), .B(dp.rf._abc_6362_n8819), .Y(dp.rf._abc_6362_n8820) );
	NAND2X1 NAND2X1_5969 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8820), .Y(dp.rf._abc_6362_n8821) );
	AND2X2 AND2X2_362 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8817), .B(dp.rf._abc_6362_n8821), .Y(dp.rf._abc_6362_n8822) );
	NAND2X1 NAND2X1_5970 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8822), .Y(dp.rf._abc_6362_n8823) );
	AND2X2 AND2X2_363 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8823), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n8824) );
	NAND2X1 NAND2X1_5971 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8813), .B(dp.rf._abc_6362_n8824), .Y(dp.rf._abc_6362_n8825) );
	NAND2X1 NAND2X1_5972 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8826) );
	NAND2X1 NAND2X1_5973 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<2>), .Y(dp.rf._abc_6362_n8827) );
	AND2X2 AND2X2_364 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8827), .B(instr[17]), .Y(dp.rf._abc_6362_n8828) );
	NAND2X1 NAND2X1_5974 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8826), .B(dp.rf._abc_6362_n8828), .Y(dp.rf._abc_6362_n8829) );
	NAND2X1 NAND2X1_5975 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8830) );
	NAND2X1 NAND2X1_5976 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<2>), .Y(dp.rf._abc_6362_n8831) );
	AND2X2 AND2X2_365 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8831), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n8832) );
	NAND2X1 NAND2X1_5977 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8830), .B(dp.rf._abc_6362_n8832), .Y(dp.rf._abc_6362_n8833) );
	NAND2X1 NAND2X1_5978 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8829), .B(dp.rf._abc_6362_n8833), .Y(dp.rf._abc_6362_n8834) );
	AND2X2 AND2X2_366 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8834), .B(instr[18]), .Y(dp.rf._abc_6362_n8835) );
	NAND2X1 NAND2X1_5979 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8836) );
	NAND2X1 NAND2X1_5980 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<2>), .Y(dp.rf._abc_6362_n8837) );
	AND2X2 AND2X2_367 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8837), .B(instr[17]), .Y(dp.rf._abc_6362_n8838) );
	NAND2X1 NAND2X1_5981 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8836), .B(dp.rf._abc_6362_n8838), .Y(dp.rf._abc_6362_n8839) );
	NAND2X1 NAND2X1_5982 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<2>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8840) );
	NAND2X1 NAND2X1_5983 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<2>), .Y(dp.rf._abc_6362_n8841) );
	AND2X2 AND2X2_368 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8841), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n8842) );
	NAND2X1 NAND2X1_5984 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8840), .B(dp.rf._abc_6362_n8842), .Y(dp.rf._abc_6362_n8843) );
	NAND2X1 NAND2X1_5985 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8839), .B(dp.rf._abc_6362_n8843), .Y(dp.rf._abc_6362_n8844) );
	NAND2X1 NAND2X1_5986 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8844), .Y(dp.rf._abc_6362_n8845) );
	NAND2X1 NAND2X1_5987 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n8845), .Y(dp.rf._abc_6362_n8846) );
	NOR2X1 NOR2X1_958 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8835), .B(dp.rf._abc_6362_n8846), .Y(dp.rf._abc_6362_n8847) );
	NOR2X1 NOR2X1_959 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n8847), .Y(dp.rf._abc_6362_n8848) );
	NAND2X1 NAND2X1_5988 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8825), .B(dp.rf._abc_6362_n8848), .Y(dp.rf._abc_6362_n8849) );
	NAND2X1 NAND2X1_5989 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n8849), .Y(dp.rf._abc_6362_n8850) );
	NOR2X1 NOR2X1_960 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8803), .B(dp.rf._abc_6362_n8850), .Y(writedata_2__RAW) );
	NAND2X1 NAND2X1_5990 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<3>), .Y(dp.rf._abc_6362_n8852) );
	NAND2X1 NAND2X1_5991 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8852), .Y(dp.rf._abc_6362_n8853) );
	NOR2X1 NOR2X1_961 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5659), .Y(dp.rf._abc_6362_n8854) );
	NOR2X1 NOR2X1_962 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8853), .B(dp.rf._abc_6362_n8854), .Y(dp.rf._abc_6362_n8855) );
	NAND2X1 NAND2X1_5992 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<3>), .Y(dp.rf._abc_6362_n8856) );
	NAND2X1 NAND2X1_5993 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8856), .Y(dp.rf._abc_6362_n8857) );
	NOR2X1 NOR2X1_963 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5664), .Y(dp.rf._abc_6362_n8858) );
	NOR2X1 NOR2X1_964 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8857), .B(dp.rf._abc_6362_n8858), .Y(dp.rf._abc_6362_n8859) );
	NOR2X1 NOR2X1_965 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8855), .B(dp.rf._abc_6362_n8859), .Y(dp.rf._abc_6362_n8860) );
	NAND2X1 NAND2X1_5994 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8860), .Y(dp.rf._abc_6362_n8861) );
	NAND2X1 NAND2X1_5995 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<3>), .Y(dp.rf._abc_6362_n8862) );
	NAND2X1 NAND2X1_5996 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8862), .Y(dp.rf._abc_6362_n8863) );
	NOR2X1 NOR2X1_966 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5671), .Y(dp.rf._abc_6362_n8864) );
	NOR2X1 NOR2X1_967 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8863), .B(dp.rf._abc_6362_n8864), .Y(dp.rf._abc_6362_n8865) );
	NAND2X1 NAND2X1_5997 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<3>), .Y(dp.rf._abc_6362_n8866) );
	NAND2X1 NAND2X1_5998 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8866), .Y(dp.rf._abc_6362_n8867) );
	NOR2X1 NOR2X1_968 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5676), .Y(dp.rf._abc_6362_n8868) );
	NOR2X1 NOR2X1_969 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8867), .B(dp.rf._abc_6362_n8868), .Y(dp.rf._abc_6362_n8869) );
	NOR2X1 NOR2X1_970 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8865), .B(dp.rf._abc_6362_n8869), .Y(dp.rf._abc_6362_n8870) );
	NAND2X1 NAND2X1_5999 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8870), .Y(dp.rf._abc_6362_n8871) );
	NAND2X1 NAND2X1_6000 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8861), .B(dp.rf._abc_6362_n8871), .Y(dp.rf._abc_6362_n8872) );
	NAND2X1 NAND2X1_6001 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n8872), .Y(dp.rf._abc_6362_n8873) );
	NAND2X1 NAND2X1_6002 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n8873), .Y(dp.rf._abc_6362_n8874) );
	NAND2X1 NAND2X1_6003 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8875) );
	NOR2X1 NOR2X1_971 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5685), .Y(dp.rf._abc_6362_n8876) );
	NOR2X1 NOR2X1_972 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8876), .Y(dp.rf._abc_6362_n8877) );
	NAND2X1 NAND2X1_6004 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8875), .B(dp.rf._abc_6362_n8877), .Y(dp.rf._abc_6362_n8878) );
	NAND2X1 NAND2X1_6005 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8879) );
	NOR2X1 NOR2X1_973 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5690), .Y(dp.rf._abc_6362_n8880) );
	NOR2X1 NOR2X1_974 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8880), .Y(dp.rf._abc_6362_n8881) );
	NAND2X1 NAND2X1_6006 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8879), .B(dp.rf._abc_6362_n8881), .Y(dp.rf._abc_6362_n8882) );
	NAND2X1 NAND2X1_6007 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8878), .B(dp.rf._abc_6362_n8882), .Y(dp.rf._abc_6362_n8883) );
	NOR2X1 NOR2X1_975 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8883), .Y(dp.rf._abc_6362_n8884) );
	NAND2X1 NAND2X1_6008 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8885) );
	NOR2X1 NOR2X1_976 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5697), .Y(dp.rf._abc_6362_n8886) );
	NOR2X1 NOR2X1_977 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8886), .Y(dp.rf._abc_6362_n8887) );
	NAND2X1 NAND2X1_6009 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8885), .B(dp.rf._abc_6362_n8887), .Y(dp.rf._abc_6362_n8888) );
	NAND2X1 NAND2X1_6010 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8889) );
	NOR2X1 NOR2X1_978 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n5702), .Y(dp.rf._abc_6362_n8890) );
	NOR2X1 NOR2X1_979 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8890), .Y(dp.rf._abc_6362_n8891) );
	NAND2X1 NAND2X1_6011 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8889), .B(dp.rf._abc_6362_n8891), .Y(dp.rf._abc_6362_n8892) );
	NAND2X1 NAND2X1_6012 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8888), .B(dp.rf._abc_6362_n8892), .Y(dp.rf._abc_6362_n8893) );
	NOR2X1 NOR2X1_980 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8893), .Y(dp.rf._abc_6362_n8894) );
	NOR2X1 NOR2X1_981 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8884), .B(dp.rf._abc_6362_n8894), .Y(dp.rf._abc_6362_n8895) );
	NOR2X1 NOR2X1_982 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n8895), .Y(dp.rf._abc_6362_n8896) );
	NOR2X1 NOR2X1_983 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8874), .B(dp.rf._abc_6362_n8896), .Y(dp.rf._abc_6362_n8897) );
	NAND2X1 NAND2X1_6013 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<3>), .Y(dp.rf._abc_6362_n8898) );
	NAND2X1 NAND2X1_6014 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8899) );
	NAND2X1 NAND2X1_6015 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8898), .B(dp.rf._abc_6362_n8899), .Y(dp.rf._abc_6362_n8900) );
	NAND2X1 NAND2X1_6016 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8900), .Y(dp.rf._abc_6362_n8901) );
	NAND2X1 NAND2X1_6017 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<3>), .Y(dp.rf._abc_6362_n8902) );
	NAND2X1 NAND2X1_6018 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8903) );
	NAND2X1 NAND2X1_6019 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8902), .B(dp.rf._abc_6362_n8903), .Y(dp.rf._abc_6362_n8904) );
	NAND2X1 NAND2X1_6020 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8904), .Y(dp.rf._abc_6362_n8905) );
	AND2X2 AND2X2_369 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8901), .B(dp.rf._abc_6362_n8905), .Y(dp.rf._abc_6362_n8906) );
	NAND2X1 NAND2X1_6021 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8906), .Y(dp.rf._abc_6362_n8907) );
	NAND2X1 NAND2X1_6022 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<3>), .Y(dp.rf._abc_6362_n8908) );
	NAND2X1 NAND2X1_6023 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8909) );
	NAND2X1 NAND2X1_6024 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8908), .B(dp.rf._abc_6362_n8909), .Y(dp.rf._abc_6362_n8910) );
	NAND2X1 NAND2X1_6025 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8910), .Y(dp.rf._abc_6362_n8911) );
	NAND2X1 NAND2X1_6026 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<3>), .Y(dp.rf._abc_6362_n8912) );
	NAND2X1 NAND2X1_6027 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8913) );
	NAND2X1 NAND2X1_6028 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8912), .B(dp.rf._abc_6362_n8913), .Y(dp.rf._abc_6362_n8914) );
	NAND2X1 NAND2X1_6029 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8914), .Y(dp.rf._abc_6362_n8915) );
	AND2X2 AND2X2_370 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8911), .B(dp.rf._abc_6362_n8915), .Y(dp.rf._abc_6362_n8916) );
	NAND2X1 NAND2X1_6030 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8916), .Y(dp.rf._abc_6362_n8917) );
	AND2X2 AND2X2_371 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8917), .B(instr[19]), .Y(dp.rf._abc_6362_n8918) );
	NAND2X1 NAND2X1_6031 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8907), .B(dp.rf._abc_6362_n8918), .Y(dp.rf._abc_6362_n8919) );
	NAND2X1 NAND2X1_6032 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8920) );
	NAND2X1 NAND2X1_6033 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<3>), .Y(dp.rf._abc_6362_n8921) );
	AND2X2 AND2X2_372 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8921), .B(instr[17]), .Y(dp.rf._abc_6362_n8922) );
	NAND2X1 NAND2X1_6034 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8920), .B(dp.rf._abc_6362_n8922), .Y(dp.rf._abc_6362_n8923) );
	NAND2X1 NAND2X1_6035 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8924) );
	NAND2X1 NAND2X1_6036 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<3>), .Y(dp.rf._abc_6362_n8925) );
	AND2X2 AND2X2_373 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8925), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n8926) );
	NAND2X1 NAND2X1_6037 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8924), .B(dp.rf._abc_6362_n8926), .Y(dp.rf._abc_6362_n8927) );
	NAND2X1 NAND2X1_6038 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8923), .B(dp.rf._abc_6362_n8927), .Y(dp.rf._abc_6362_n8928) );
	AND2X2 AND2X2_374 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8928), .B(instr[18]), .Y(dp.rf._abc_6362_n8929) );
	NAND2X1 NAND2X1_6039 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8930) );
	NAND2X1 NAND2X1_6040 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<3>), .Y(dp.rf._abc_6362_n8931) );
	AND2X2 AND2X2_375 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8931), .B(instr[17]), .Y(dp.rf._abc_6362_n8932) );
	NAND2X1 NAND2X1_6041 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8930), .B(dp.rf._abc_6362_n8932), .Y(dp.rf._abc_6362_n8933) );
	NAND2X1 NAND2X1_6042 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<3>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8934) );
	NAND2X1 NAND2X1_6043 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<3>), .Y(dp.rf._abc_6362_n8935) );
	AND2X2 AND2X2_376 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8935), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n8936) );
	NAND2X1 NAND2X1_6044 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8934), .B(dp.rf._abc_6362_n8936), .Y(dp.rf._abc_6362_n8937) );
	NAND2X1 NAND2X1_6045 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8933), .B(dp.rf._abc_6362_n8937), .Y(dp.rf._abc_6362_n8938) );
	NAND2X1 NAND2X1_6046 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8938), .Y(dp.rf._abc_6362_n8939) );
	NAND2X1 NAND2X1_6047 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n8939), .Y(dp.rf._abc_6362_n8940) );
	NOR2X1 NOR2X1_984 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8929), .B(dp.rf._abc_6362_n8940), .Y(dp.rf._abc_6362_n8941) );
	NOR2X1 NOR2X1_985 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n8941), .Y(dp.rf._abc_6362_n8942) );
	NAND2X1 NAND2X1_6048 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8919), .B(dp.rf._abc_6362_n8942), .Y(dp.rf._abc_6362_n8943) );
	NAND2X1 NAND2X1_6049 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n8943), .Y(dp.rf._abc_6362_n8944) );
	NOR2X1 NOR2X1_986 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8897), .B(dp.rf._abc_6362_n8944), .Y(writedata_3__RAW) );
	NAND2X1 NAND2X1_6050 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<4>), .Y(dp.rf._abc_6362_n8946) );
	NAND2X1 NAND2X1_6051 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8946), .Y(dp.rf._abc_6362_n8947) );
	NOR2X1 NOR2X1_987 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5783), .Y(dp.rf._abc_6362_n8948) );
	NOR2X1 NOR2X1_988 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8947), .B(dp.rf._abc_6362_n8948), .Y(dp.rf._abc_6362_n8949) );
	NAND2X1 NAND2X1_6052 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<4>), .Y(dp.rf._abc_6362_n8950) );
	NAND2X1 NAND2X1_6053 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8950), .Y(dp.rf._abc_6362_n8951) );
	NOR2X1 NOR2X1_989 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5788), .Y(dp.rf._abc_6362_n8952) );
	NOR2X1 NOR2X1_990 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8951), .B(dp.rf._abc_6362_n8952), .Y(dp.rf._abc_6362_n8953) );
	NOR2X1 NOR2X1_991 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8949), .B(dp.rf._abc_6362_n8953), .Y(dp.rf._abc_6362_n8954) );
	NAND2X1 NAND2X1_6054 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8954), .Y(dp.rf._abc_6362_n8955) );
	NAND2X1 NAND2X1_6055 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<4>), .Y(dp.rf._abc_6362_n8956) );
	NAND2X1 NAND2X1_6056 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8956), .Y(dp.rf._abc_6362_n8957) );
	NOR2X1 NOR2X1_992 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5795), .Y(dp.rf._abc_6362_n8958) );
	NOR2X1 NOR2X1_993 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8957), .B(dp.rf._abc_6362_n8958), .Y(dp.rf._abc_6362_n8959) );
	NAND2X1 NAND2X1_6057 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<4>), .Y(dp.rf._abc_6362_n8960) );
	NAND2X1 NAND2X1_6058 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8960), .Y(dp.rf._abc_6362_n8961) );
	NOR2X1 NOR2X1_994 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5800), .Y(dp.rf._abc_6362_n8962) );
	NOR2X1 NOR2X1_995 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8961), .B(dp.rf._abc_6362_n8962), .Y(dp.rf._abc_6362_n8963) );
	NOR2X1 NOR2X1_996 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8959), .B(dp.rf._abc_6362_n8963), .Y(dp.rf._abc_6362_n8964) );
	NAND2X1 NAND2X1_6059 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8964), .Y(dp.rf._abc_6362_n8965) );
	NAND2X1 NAND2X1_6060 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8955), .B(dp.rf._abc_6362_n8965), .Y(dp.rf._abc_6362_n8966) );
	NAND2X1 NAND2X1_6061 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n8966), .Y(dp.rf._abc_6362_n8967) );
	NAND2X1 NAND2X1_6062 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<4>), .Y(dp.rf._abc_6362_n8968) );
	NAND2X1 NAND2X1_6063 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<4>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8969) );
	NAND2X1 NAND2X1_6064 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8968), .B(dp.rf._abc_6362_n8969), .Y(dp.rf._abc_6362_n8970) );
	NAND2X1 NAND2X1_6065 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8970), .Y(dp.rf._abc_6362_n8971) );
	NAND2X1 NAND2X1_6066 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<4>), .Y(dp.rf._abc_6362_n8972) );
	NAND2X1 NAND2X1_6067 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<4>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8973) );
	NAND2X1 NAND2X1_6068 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8972), .B(dp.rf._abc_6362_n8973), .Y(dp.rf._abc_6362_n8974) );
	NAND2X1 NAND2X1_6069 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8974), .Y(dp.rf._abc_6362_n8975) );
	AND2X2 AND2X2_377 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8971), .B(dp.rf._abc_6362_n8975), .Y(dp.rf._abc_6362_n8976) );
	NAND2X1 NAND2X1_6070 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n8976), .Y(dp.rf._abc_6362_n8977) );
	NAND2X1 NAND2X1_6071 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<4>), .Y(dp.rf._abc_6362_n8978) );
	NAND2X1 NAND2X1_6072 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8978), .Y(dp.rf._abc_6362_n8979) );
	AND2X2 AND2X2_378 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf.rf_2_<4>), .Y(dp.rf._abc_6362_n8980) );
	NOR2X1 NOR2X1_997 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8979), .B(dp.rf._abc_6362_n8980), .Y(dp.rf._abc_6362_n8981) );
	NAND2X1 NAND2X1_6073 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<4>), .Y(dp.rf._abc_6362_n8982) );
	NAND2X1 NAND2X1_6074 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8982), .Y(dp.rf._abc_6362_n8983) );
	INVX1 INVX1_254 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<4>), .Y(dp.rf._abc_6362_n8984) );
	NOR2X1 NOR2X1_998 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8984), .Y(dp.rf._abc_6362_n8985) );
	NOR2X1 NOR2X1_999 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8983), .B(dp.rf._abc_6362_n8985), .Y(dp.rf._abc_6362_n8986) );
	OR2X2 OR2X2_86 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8981), .B(dp.rf._abc_6362_n8986), .Y(dp.rf._abc_6362_n8987) );
	NAND2X1 NAND2X1_6075 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n8987), .Y(dp.rf._abc_6362_n8988) );
	AND2X2 AND2X2_379 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8988), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n8989) );
	NAND2X1 NAND2X1_6076 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8977), .B(dp.rf._abc_6362_n8989), .Y(dp.rf._abc_6362_n8990) );
	NAND2X1 NAND2X1_6077 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8967), .B(dp.rf._abc_6362_n8990), .Y(dp.rf._abc_6362_n8991) );
	NOR2X1 NOR2X1_1000 ( .gnd(gnd), .vdd(vdd), .A(instr[20]), .B(dp.rf._abc_6362_n8991), .Y(dp.rf._abc_6362_n8992) );
	NAND2X1 NAND2X1_6078 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<4>), .Y(dp.rf._abc_6362_n8993) );
	NAND2X1 NAND2X1_6079 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<4>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8994) );
	NAND2X1 NAND2X1_6080 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8993), .B(dp.rf._abc_6362_n8994), .Y(dp.rf._abc_6362_n8995) );
	NAND2X1 NAND2X1_6081 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n8995), .Y(dp.rf._abc_6362_n8996) );
	NAND2X1 NAND2X1_6082 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<4>), .Y(dp.rf._abc_6362_n8997) );
	NAND2X1 NAND2X1_6083 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<4>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n8998) );
	NAND2X1 NAND2X1_6084 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8997), .B(dp.rf._abc_6362_n8998), .Y(dp.rf._abc_6362_n8999) );
	NAND2X1 NAND2X1_6085 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n8999), .Y(dp.rf._abc_6362_n9000) );
	AND2X2 AND2X2_380 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8996), .B(dp.rf._abc_6362_n9000), .Y(dp.rf._abc_6362_n9001) );
	NAND2X1 NAND2X1_6086 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9001), .Y(dp.rf._abc_6362_n9002) );
	NAND2X1 NAND2X1_6087 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<4>), .Y(dp.rf._abc_6362_n9003) );
	NAND2X1 NAND2X1_6088 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<4>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9004) );
	NAND2X1 NAND2X1_6089 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9003), .B(dp.rf._abc_6362_n9004), .Y(dp.rf._abc_6362_n9005) );
	NAND2X1 NAND2X1_6090 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9005), .Y(dp.rf._abc_6362_n9006) );
	NAND2X1 NAND2X1_6091 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<4>), .Y(dp.rf._abc_6362_n9007) );
	NAND2X1 NAND2X1_6092 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<4>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9008) );
	NAND2X1 NAND2X1_6093 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9007), .B(dp.rf._abc_6362_n9008), .Y(dp.rf._abc_6362_n9009) );
	NAND2X1 NAND2X1_6094 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9009), .Y(dp.rf._abc_6362_n9010) );
	AND2X2 AND2X2_381 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9006), .B(dp.rf._abc_6362_n9010), .Y(dp.rf._abc_6362_n9011) );
	NAND2X1 NAND2X1_6095 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9011), .Y(dp.rf._abc_6362_n9012) );
	AND2X2 AND2X2_382 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9012), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n9013) );
	NAND2X1 NAND2X1_6096 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9002), .B(dp.rf._abc_6362_n9013), .Y(dp.rf._abc_6362_n9014) );
	NAND2X1 NAND2X1_6097 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<4>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9015) );
	NAND2X1 NAND2X1_6098 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<4>), .Y(dp.rf._abc_6362_n9016) );
	AND2X2 AND2X2_383 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9016), .B(instr[17]), .Y(dp.rf._abc_6362_n9017) );
	NAND2X1 NAND2X1_6099 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9015), .B(dp.rf._abc_6362_n9017), .Y(dp.rf._abc_6362_n9018) );
	NAND2X1 NAND2X1_6100 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<4>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9019) );
	NAND2X1 NAND2X1_6101 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<4>), .Y(dp.rf._abc_6362_n9020) );
	AND2X2 AND2X2_384 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9020), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9021) );
	NAND2X1 NAND2X1_6102 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9019), .B(dp.rf._abc_6362_n9021), .Y(dp.rf._abc_6362_n9022) );
	NAND2X1 NAND2X1_6103 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9018), .B(dp.rf._abc_6362_n9022), .Y(dp.rf._abc_6362_n9023) );
	AND2X2 AND2X2_385 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9023), .B(instr[18]), .Y(dp.rf._abc_6362_n9024) );
	NAND2X1 NAND2X1_6104 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<4>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9025) );
	NAND2X1 NAND2X1_6105 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<4>), .Y(dp.rf._abc_6362_n9026) );
	AND2X2 AND2X2_386 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9026), .B(instr[17]), .Y(dp.rf._abc_6362_n9027) );
	NAND2X1 NAND2X1_6106 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9025), .B(dp.rf._abc_6362_n9027), .Y(dp.rf._abc_6362_n9028) );
	NAND2X1 NAND2X1_6107 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<4>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9029) );
	NAND2X1 NAND2X1_6108 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<4>), .Y(dp.rf._abc_6362_n9030) );
	AND2X2 AND2X2_387 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9030), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9031) );
	NAND2X1 NAND2X1_6109 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9029), .B(dp.rf._abc_6362_n9031), .Y(dp.rf._abc_6362_n9032) );
	NAND2X1 NAND2X1_6110 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9028), .B(dp.rf._abc_6362_n9032), .Y(dp.rf._abc_6362_n9033) );
	NAND2X1 NAND2X1_6111 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9033), .Y(dp.rf._abc_6362_n9034) );
	NAND2X1 NAND2X1_6112 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9034), .Y(dp.rf._abc_6362_n9035) );
	NOR2X1 NOR2X1_1001 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9024), .B(dp.rf._abc_6362_n9035), .Y(dp.rf._abc_6362_n9036) );
	NOR2X1 NOR2X1_1002 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9036), .Y(dp.rf._abc_6362_n9037) );
	NAND2X1 NAND2X1_6113 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9014), .B(dp.rf._abc_6362_n9037), .Y(dp.rf._abc_6362_n9038) );
	NAND2X1 NAND2X1_6114 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n9038), .Y(dp.rf._abc_6362_n9039) );
	NOR2X1 NOR2X1_1003 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8992), .B(dp.rf._abc_6362_n9039), .Y(writedata_4__RAW) );
	NAND2X1 NAND2X1_6115 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<5>), .Y(dp.rf._abc_6362_n9041) );
	NAND2X1 NAND2X1_6116 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9042) );
	NAND2X1 NAND2X1_6117 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9041), .B(dp.rf._abc_6362_n9042), .Y(dp.rf._abc_6362_n9043) );
	NAND2X1 NAND2X1_6118 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9043), .Y(dp.rf._abc_6362_n9044) );
	NAND2X1 NAND2X1_6119 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<5>), .Y(dp.rf._abc_6362_n9045) );
	NAND2X1 NAND2X1_6120 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9046) );
	NAND2X1 NAND2X1_6121 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9045), .B(dp.rf._abc_6362_n9046), .Y(dp.rf._abc_6362_n9047) );
	NAND2X1 NAND2X1_6122 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9047), .Y(dp.rf._abc_6362_n9048) );
	NAND2X1 NAND2X1_6123 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9044), .B(dp.rf._abc_6362_n9048), .Y(dp.rf._abc_6362_n9049) );
	NOR2X1 NOR2X1_1004 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9049), .Y(dp.rf._abc_6362_n9050) );
	NAND2X1 NAND2X1_6124 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<5>), .Y(dp.rf._abc_6362_n9051) );
	NAND2X1 NAND2X1_6125 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9052) );
	NAND2X1 NAND2X1_6126 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9051), .B(dp.rf._abc_6362_n9052), .Y(dp.rf._abc_6362_n9053) );
	NAND2X1 NAND2X1_6127 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9053), .Y(dp.rf._abc_6362_n9054) );
	NAND2X1 NAND2X1_6128 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<5>), .Y(dp.rf._abc_6362_n9055) );
	NAND2X1 NAND2X1_6129 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9056) );
	NAND2X1 NAND2X1_6130 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9055), .B(dp.rf._abc_6362_n9056), .Y(dp.rf._abc_6362_n9057) );
	NAND2X1 NAND2X1_6131 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9057), .Y(dp.rf._abc_6362_n9058) );
	AND2X2 AND2X2_388 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9054), .B(dp.rf._abc_6362_n9058), .Y(dp.rf._abc_6362_n9059) );
	NAND2X1 NAND2X1_6132 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9059), .Y(dp.rf._abc_6362_n9060) );
	NAND2X1 NAND2X1_6133 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n9060), .Y(dp.rf._abc_6362_n9061) );
	NOR2X1 NOR2X1_1005 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9050), .B(dp.rf._abc_6362_n9061), .Y(dp.rf._abc_6362_n9062) );
	NAND2X1 NAND2X1_6134 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<5>), .Y(dp.rf._abc_6362_n9063) );
	NAND2X1 NAND2X1_6135 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9064) );
	NAND2X1 NAND2X1_6136 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9063), .B(dp.rf._abc_6362_n9064), .Y(dp.rf._abc_6362_n9065) );
	NAND2X1 NAND2X1_6137 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9065), .Y(dp.rf._abc_6362_n9066) );
	NAND2X1 NAND2X1_6138 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<5>), .Y(dp.rf._abc_6362_n9067) );
	NAND2X1 NAND2X1_6139 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9068) );
	NAND2X1 NAND2X1_6140 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9067), .B(dp.rf._abc_6362_n9068), .Y(dp.rf._abc_6362_n9069) );
	NAND2X1 NAND2X1_6141 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9069), .Y(dp.rf._abc_6362_n9070) );
	NAND2X1 NAND2X1_6142 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9066), .B(dp.rf._abc_6362_n9070), .Y(dp.rf._abc_6362_n9071) );
	NAND2X1 NAND2X1_6143 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9071), .Y(dp.rf._abc_6362_n9072) );
	NAND2X1 NAND2X1_6144 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<5>), .Y(dp.rf._abc_6362_n9073) );
	NAND2X1 NAND2X1_6145 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9074) );
	NAND2X1 NAND2X1_6146 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9073), .B(dp.rf._abc_6362_n9074), .Y(dp.rf._abc_6362_n9075) );
	NAND2X1 NAND2X1_6147 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9075), .Y(dp.rf._abc_6362_n9076) );
	NAND2X1 NAND2X1_6148 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<5>), .Y(dp.rf._abc_6362_n9077) );
	NAND2X1 NAND2X1_6149 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9078) );
	NAND2X1 NAND2X1_6150 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9077), .B(dp.rf._abc_6362_n9078), .Y(dp.rf._abc_6362_n9079) );
	NAND2X1 NAND2X1_6151 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9079), .Y(dp.rf._abc_6362_n9080) );
	NAND2X1 NAND2X1_6152 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9076), .B(dp.rf._abc_6362_n9080), .Y(dp.rf._abc_6362_n9081) );
	NAND2X1 NAND2X1_6153 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9081), .Y(dp.rf._abc_6362_n9082) );
	NAND2X1 NAND2X1_6154 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9072), .B(dp.rf._abc_6362_n9082), .Y(dp.rf._abc_6362_n9083) );
	NAND2X1 NAND2X1_6155 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9083), .Y(dp.rf._abc_6362_n9084) );
	NAND2X1 NAND2X1_6156 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9084), .Y(dp.rf._abc_6362_n9085) );
	NOR2X1 NOR2X1_1006 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9062), .B(dp.rf._abc_6362_n9085), .Y(dp.rf._abc_6362_n9086) );
	NAND2X1 NAND2X1_6157 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<5>), .Y(dp.rf._abc_6362_n9087) );
	NAND2X1 NAND2X1_6158 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9087), .Y(dp.rf._abc_6362_n9088) );
	NOR2X1 NOR2X1_1007 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5906), .Y(dp.rf._abc_6362_n9089) );
	NOR2X1 NOR2X1_1008 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9088), .B(dp.rf._abc_6362_n9089), .Y(dp.rf._abc_6362_n9090) );
	NAND2X1 NAND2X1_6159 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<5>), .Y(dp.rf._abc_6362_n9091) );
	NAND2X1 NAND2X1_6160 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9091), .Y(dp.rf._abc_6362_n9092) );
	NOR2X1 NOR2X1_1009 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5911), .Y(dp.rf._abc_6362_n9093) );
	NOR2X1 NOR2X1_1010 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9092), .B(dp.rf._abc_6362_n9093), .Y(dp.rf._abc_6362_n9094) );
	OR2X2 OR2X2_87 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9090), .B(dp.rf._abc_6362_n9094), .Y(dp.rf._abc_6362_n9095) );
	NAND2X1 NAND2X1_6161 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9095), .Y(dp.rf._abc_6362_n9096) );
	NAND2X1 NAND2X1_6162 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<5>), .Y(dp.rf._abc_6362_n9097) );
	NAND2X1 NAND2X1_6163 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9097), .Y(dp.rf._abc_6362_n9098) );
	NOR2X1 NOR2X1_1011 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5918), .Y(dp.rf._abc_6362_n9099) );
	NOR2X1 NOR2X1_1012 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9098), .B(dp.rf._abc_6362_n9099), .Y(dp.rf._abc_6362_n9100) );
	NAND2X1 NAND2X1_6164 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<5>), .Y(dp.rf._abc_6362_n9101) );
	NAND2X1 NAND2X1_6165 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9101), .Y(dp.rf._abc_6362_n9102) );
	NOR2X1 NOR2X1_1013 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n5923), .Y(dp.rf._abc_6362_n9103) );
	NOR2X1 NOR2X1_1014 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9102), .B(dp.rf._abc_6362_n9103), .Y(dp.rf._abc_6362_n9104) );
	OR2X2 OR2X2_88 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9100), .B(dp.rf._abc_6362_n9104), .Y(dp.rf._abc_6362_n9105) );
	NAND2X1 NAND2X1_6166 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9105), .Y(dp.rf._abc_6362_n9106) );
	AND2X2 AND2X2_389 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9106), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n9107) );
	NAND2X1 NAND2X1_6167 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9096), .B(dp.rf._abc_6362_n9107), .Y(dp.rf._abc_6362_n9108) );
	NAND2X1 NAND2X1_6168 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9109) );
	NAND2X1 NAND2X1_6169 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<5>), .Y(dp.rf._abc_6362_n9110) );
	AND2X2 AND2X2_390 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9110), .B(instr[17]), .Y(dp.rf._abc_6362_n9111) );
	NAND2X1 NAND2X1_6170 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9109), .B(dp.rf._abc_6362_n9111), .Y(dp.rf._abc_6362_n9112) );
	NAND2X1 NAND2X1_6171 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9113) );
	NAND2X1 NAND2X1_6172 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<5>), .Y(dp.rf._abc_6362_n9114) );
	AND2X2 AND2X2_391 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9114), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9115) );
	NAND2X1 NAND2X1_6173 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9113), .B(dp.rf._abc_6362_n9115), .Y(dp.rf._abc_6362_n9116) );
	NAND2X1 NAND2X1_6174 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9112), .B(dp.rf._abc_6362_n9116), .Y(dp.rf._abc_6362_n9117) );
	AND2X2 AND2X2_392 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9117), .B(instr[18]), .Y(dp.rf._abc_6362_n9118) );
	NAND2X1 NAND2X1_6175 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9119) );
	NAND2X1 NAND2X1_6176 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<5>), .Y(dp.rf._abc_6362_n9120) );
	AND2X2 AND2X2_393 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9120), .B(instr[17]), .Y(dp.rf._abc_6362_n9121) );
	NAND2X1 NAND2X1_6177 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9119), .B(dp.rf._abc_6362_n9121), .Y(dp.rf._abc_6362_n9122) );
	NAND2X1 NAND2X1_6178 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<5>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9123) );
	NAND2X1 NAND2X1_6179 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<5>), .Y(dp.rf._abc_6362_n9124) );
	AND2X2 AND2X2_394 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9124), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9125) );
	NAND2X1 NAND2X1_6180 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9123), .B(dp.rf._abc_6362_n9125), .Y(dp.rf._abc_6362_n9126) );
	NAND2X1 NAND2X1_6181 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9122), .B(dp.rf._abc_6362_n9126), .Y(dp.rf._abc_6362_n9127) );
	NAND2X1 NAND2X1_6182 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9127), .Y(dp.rf._abc_6362_n9128) );
	NAND2X1 NAND2X1_6183 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9128), .Y(dp.rf._abc_6362_n9129) );
	NOR2X1 NOR2X1_1015 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9118), .B(dp.rf._abc_6362_n9129), .Y(dp.rf._abc_6362_n9130) );
	NOR2X1 NOR2X1_1016 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9130), .Y(dp.rf._abc_6362_n9131) );
	NAND2X1 NAND2X1_6184 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9108), .B(dp.rf._abc_6362_n9131), .Y(dp.rf._abc_6362_n9132) );
	NAND2X1 NAND2X1_6185 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n9132), .Y(dp.rf._abc_6362_n9133) );
	NOR2X1 NOR2X1_1017 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9086), .B(dp.rf._abc_6362_n9133), .Y(writedata_5__RAW) );
	NAND2X1 NAND2X1_6186 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<6>), .Y(dp.rf._abc_6362_n9135) );
	NAND2X1 NAND2X1_6187 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<6>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9136) );
	NAND2X1 NAND2X1_6188 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9135), .B(dp.rf._abc_6362_n9136), .Y(dp.rf._abc_6362_n9137) );
	NAND2X1 NAND2X1_6189 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9137), .Y(dp.rf._abc_6362_n9138) );
	NAND2X1 NAND2X1_6190 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<6>), .Y(dp.rf._abc_6362_n9139) );
	NAND2X1 NAND2X1_6191 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<6>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9140) );
	NAND2X1 NAND2X1_6192 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9139), .B(dp.rf._abc_6362_n9140), .Y(dp.rf._abc_6362_n9141) );
	NAND2X1 NAND2X1_6193 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9141), .Y(dp.rf._abc_6362_n9142) );
	NAND2X1 NAND2X1_6194 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9138), .B(dp.rf._abc_6362_n9142), .Y(dp.rf._abc_6362_n9143) );
	NOR2X1 NOR2X1_1018 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9143), .Y(dp.rf._abc_6362_n9144) );
	NAND2X1 NAND2X1_6195 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<6>), .Y(dp.rf._abc_6362_n9145) );
	NAND2X1 NAND2X1_6196 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<6>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9146) );
	NAND2X1 NAND2X1_6197 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9145), .B(dp.rf._abc_6362_n9146), .Y(dp.rf._abc_6362_n9147) );
	NAND2X1 NAND2X1_6198 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9147), .Y(dp.rf._abc_6362_n9148) );
	NAND2X1 NAND2X1_6199 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<6>), .Y(dp.rf._abc_6362_n9149) );
	NAND2X1 NAND2X1_6200 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<6>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9150) );
	NAND2X1 NAND2X1_6201 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9149), .B(dp.rf._abc_6362_n9150), .Y(dp.rf._abc_6362_n9151) );
	NAND2X1 NAND2X1_6202 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9151), .Y(dp.rf._abc_6362_n9152) );
	AND2X2 AND2X2_395 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9148), .B(dp.rf._abc_6362_n9152), .Y(dp.rf._abc_6362_n9153) );
	NAND2X1 NAND2X1_6203 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9153), .Y(dp.rf._abc_6362_n9154) );
	NAND2X1 NAND2X1_6204 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9154), .Y(dp.rf._abc_6362_n9155) );
	NOR2X1 NOR2X1_1019 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9144), .B(dp.rf._abc_6362_n9155), .Y(dp.rf._abc_6362_n9156) );
	NAND2X1 NAND2X1_6205 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<6>), .Y(dp.rf._abc_6362_n9157) );
	NAND2X1 NAND2X1_6206 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<6>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9158) );
	NAND2X1 NAND2X1_6207 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9157), .B(dp.rf._abc_6362_n9158), .Y(dp.rf._abc_6362_n9159) );
	NAND2X1 NAND2X1_6208 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9159), .Y(dp.rf._abc_6362_n9160) );
	NAND2X1 NAND2X1_6209 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<6>), .Y(dp.rf._abc_6362_n9161) );
	NAND2X1 NAND2X1_6210 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<6>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9162) );
	NAND2X1 NAND2X1_6211 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9161), .B(dp.rf._abc_6362_n9162), .Y(dp.rf._abc_6362_n9163) );
	NAND2X1 NAND2X1_6212 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9163), .Y(dp.rf._abc_6362_n9164) );
	AND2X2 AND2X2_396 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9160), .B(dp.rf._abc_6362_n9164), .Y(dp.rf._abc_6362_n9165) );
	NAND2X1 NAND2X1_6213 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9165), .Y(dp.rf._abc_6362_n9166) );
	NAND2X1 NAND2X1_6214 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<6>), .Y(dp.rf._abc_6362_n9167) );
	NAND2X1 NAND2X1_6215 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9167), .Y(dp.rf._abc_6362_n9168) );
	AND2X2 AND2X2_397 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf.rf_2_<6>), .Y(dp.rf._abc_6362_n9169) );
	NOR2X1 NOR2X1_1020 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9168), .B(dp.rf._abc_6362_n9169), .Y(dp.rf._abc_6362_n9170) );
	NAND2X1 NAND2X1_6216 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<6>), .Y(dp.rf._abc_6362_n9171) );
	NAND2X1 NAND2X1_6217 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9171), .Y(dp.rf._abc_6362_n9172) );
	INVX1 INVX1_255 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<6>), .Y(dp.rf._abc_6362_n9173) );
	NOR2X1 NOR2X1_1021 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n9173), .Y(dp.rf._abc_6362_n9174) );
	NOR2X1 NOR2X1_1022 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9172), .B(dp.rf._abc_6362_n9174), .Y(dp.rf._abc_6362_n9175) );
	OR2X2 OR2X2_89 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9170), .B(dp.rf._abc_6362_n9175), .Y(dp.rf._abc_6362_n9176) );
	NAND2X1 NAND2X1_6218 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9176), .Y(dp.rf._abc_6362_n9177) );
	AND2X2 AND2X2_398 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9177), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n9178) );
	NAND2X1 NAND2X1_6219 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9166), .B(dp.rf._abc_6362_n9178), .Y(dp.rf._abc_6362_n9179) );
	NAND2X1 NAND2X1_6220 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9179), .Y(dp.rf._abc_6362_n9180) );
	NOR2X1 NOR2X1_1023 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9156), .B(dp.rf._abc_6362_n9180), .Y(dp.rf._abc_6362_n9181) );
	NAND2X1 NAND2X1_6221 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<6>), .Y(dp.rf._abc_6362_n9182) );
	NAND2X1 NAND2X1_6222 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9182), .Y(dp.rf._abc_6362_n9183) );
	NOR2X1 NOR2X1_1024 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6004), .Y(dp.rf._abc_6362_n9184) );
	NOR2X1 NOR2X1_1025 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9183), .B(dp.rf._abc_6362_n9184), .Y(dp.rf._abc_6362_n9185) );
	NAND2X1 NAND2X1_6223 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<6>), .Y(dp.rf._abc_6362_n9186) );
	NAND2X1 NAND2X1_6224 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9186), .Y(dp.rf._abc_6362_n9187) );
	NOR2X1 NOR2X1_1026 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6009), .Y(dp.rf._abc_6362_n9188) );
	NOR2X1 NOR2X1_1027 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9187), .B(dp.rf._abc_6362_n9188), .Y(dp.rf._abc_6362_n9189) );
	OR2X2 OR2X2_90 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9185), .B(dp.rf._abc_6362_n9189), .Y(dp.rf._abc_6362_n9190) );
	NAND2X1 NAND2X1_6225 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9190), .Y(dp.rf._abc_6362_n9191) );
	NAND2X1 NAND2X1_6226 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<6>), .Y(dp.rf._abc_6362_n9192) );
	NAND2X1 NAND2X1_6227 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9192), .Y(dp.rf._abc_6362_n9193) );
	NOR2X1 NOR2X1_1028 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6016), .Y(dp.rf._abc_6362_n9194) );
	NOR2X1 NOR2X1_1029 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9193), .B(dp.rf._abc_6362_n9194), .Y(dp.rf._abc_6362_n9195) );
	NAND2X1 NAND2X1_6228 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<6>), .Y(dp.rf._abc_6362_n9196) );
	NAND2X1 NAND2X1_6229 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9196), .Y(dp.rf._abc_6362_n9197) );
	NOR2X1 NOR2X1_1030 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6021), .Y(dp.rf._abc_6362_n9198) );
	NOR2X1 NOR2X1_1031 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9197), .B(dp.rf._abc_6362_n9198), .Y(dp.rf._abc_6362_n9199) );
	OR2X2 OR2X2_91 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9195), .B(dp.rf._abc_6362_n9199), .Y(dp.rf._abc_6362_n9200) );
	NAND2X1 NAND2X1_6230 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9200), .Y(dp.rf._abc_6362_n9201) );
	AND2X2 AND2X2_399 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9201), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n9202) );
	NAND2X1 NAND2X1_6231 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9191), .B(dp.rf._abc_6362_n9202), .Y(dp.rf._abc_6362_n9203) );
	NAND2X1 NAND2X1_6232 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<6>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9204) );
	NAND2X1 NAND2X1_6233 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<6>), .Y(dp.rf._abc_6362_n9205) );
	AND2X2 AND2X2_400 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9205), .B(instr[17]), .Y(dp.rf._abc_6362_n9206) );
	NAND2X1 NAND2X1_6234 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9204), .B(dp.rf._abc_6362_n9206), .Y(dp.rf._abc_6362_n9207) );
	NAND2X1 NAND2X1_6235 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<6>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9208) );
	NAND2X1 NAND2X1_6236 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<6>), .Y(dp.rf._abc_6362_n9209) );
	AND2X2 AND2X2_401 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9209), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9210) );
	NAND2X1 NAND2X1_6237 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9208), .B(dp.rf._abc_6362_n9210), .Y(dp.rf._abc_6362_n9211) );
	NAND2X1 NAND2X1_6238 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9207), .B(dp.rf._abc_6362_n9211), .Y(dp.rf._abc_6362_n9212) );
	AND2X2 AND2X2_402 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9212), .B(instr[18]), .Y(dp.rf._abc_6362_n9213) );
	NAND2X1 NAND2X1_6239 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<6>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9214) );
	NAND2X1 NAND2X1_6240 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<6>), .Y(dp.rf._abc_6362_n9215) );
	AND2X2 AND2X2_403 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9215), .B(instr[17]), .Y(dp.rf._abc_6362_n9216) );
	NAND2X1 NAND2X1_6241 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9214), .B(dp.rf._abc_6362_n9216), .Y(dp.rf._abc_6362_n9217) );
	NAND2X1 NAND2X1_6242 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<6>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9218) );
	NAND2X1 NAND2X1_6243 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<6>), .Y(dp.rf._abc_6362_n9219) );
	AND2X2 AND2X2_404 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9219), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9220) );
	NAND2X1 NAND2X1_6244 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9218), .B(dp.rf._abc_6362_n9220), .Y(dp.rf._abc_6362_n9221) );
	NAND2X1 NAND2X1_6245 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9217), .B(dp.rf._abc_6362_n9221), .Y(dp.rf._abc_6362_n9222) );
	NAND2X1 NAND2X1_6246 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9222), .Y(dp.rf._abc_6362_n9223) );
	NAND2X1 NAND2X1_6247 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9223), .Y(dp.rf._abc_6362_n9224) );
	NOR2X1 NOR2X1_1032 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9213), .B(dp.rf._abc_6362_n9224), .Y(dp.rf._abc_6362_n9225) );
	NOR2X1 NOR2X1_1033 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9225), .Y(dp.rf._abc_6362_n9226) );
	NAND2X1 NAND2X1_6248 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9203), .B(dp.rf._abc_6362_n9226), .Y(dp.rf._abc_6362_n9227) );
	NAND2X1 NAND2X1_6249 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n9227), .Y(dp.rf._abc_6362_n9228) );
	NOR2X1 NOR2X1_1034 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9181), .B(dp.rf._abc_6362_n9228), .Y(writedata_6__RAW) );
	NAND2X1 NAND2X1_6250 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<7>), .Y(dp.rf._abc_6362_n9230) );
	NAND2X1 NAND2X1_6251 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<7>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9231) );
	NAND2X1 NAND2X1_6252 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9230), .B(dp.rf._abc_6362_n9231), .Y(dp.rf._abc_6362_n9232) );
	NAND2X1 NAND2X1_6253 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9232), .Y(dp.rf._abc_6362_n9233) );
	NAND2X1 NAND2X1_6254 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<7>), .Y(dp.rf._abc_6362_n9234) );
	NAND2X1 NAND2X1_6255 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<7>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9235) );
	NAND2X1 NAND2X1_6256 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9234), .B(dp.rf._abc_6362_n9235), .Y(dp.rf._abc_6362_n9236) );
	NAND2X1 NAND2X1_6257 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9236), .Y(dp.rf._abc_6362_n9237) );
	NAND2X1 NAND2X1_6258 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9233), .B(dp.rf._abc_6362_n9237), .Y(dp.rf._abc_6362_n9238) );
	NOR2X1 NOR2X1_1035 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9238), .Y(dp.rf._abc_6362_n9239) );
	NAND2X1 NAND2X1_6259 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<7>), .Y(dp.rf._abc_6362_n9240) );
	NAND2X1 NAND2X1_6260 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<7>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9241) );
	NAND2X1 NAND2X1_6261 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9240), .B(dp.rf._abc_6362_n9241), .Y(dp.rf._abc_6362_n9242) );
	NAND2X1 NAND2X1_6262 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9242), .Y(dp.rf._abc_6362_n9243) );
	NAND2X1 NAND2X1_6263 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<7>), .Y(dp.rf._abc_6362_n9244) );
	NAND2X1 NAND2X1_6264 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<7>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9245) );
	NAND2X1 NAND2X1_6265 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9244), .B(dp.rf._abc_6362_n9245), .Y(dp.rf._abc_6362_n9246) );
	NAND2X1 NAND2X1_6266 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9246), .Y(dp.rf._abc_6362_n9247) );
	AND2X2 AND2X2_405 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9243), .B(dp.rf._abc_6362_n9247), .Y(dp.rf._abc_6362_n9248) );
	NAND2X1 NAND2X1_6267 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9248), .Y(dp.rf._abc_6362_n9249) );
	NAND2X1 NAND2X1_6268 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n9249), .Y(dp.rf._abc_6362_n9250) );
	NOR2X1 NOR2X1_1036 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9239), .B(dp.rf._abc_6362_n9250), .Y(dp.rf._abc_6362_n9251) );
	NAND2X1 NAND2X1_6269 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<7>), .Y(dp.rf._abc_6362_n9252) );
	NAND2X1 NAND2X1_6270 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9252), .Y(dp.rf._abc_6362_n9253) );
	NOR2X1 NOR2X1_1037 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6056), .Y(dp.rf._abc_6362_n9254) );
	NOR2X1 NOR2X1_1038 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9253), .B(dp.rf._abc_6362_n9254), .Y(dp.rf._abc_6362_n9255) );
	NAND2X1 NAND2X1_6271 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<7>), .Y(dp.rf._abc_6362_n9256) );
	NAND2X1 NAND2X1_6272 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9256), .Y(dp.rf._abc_6362_n9257) );
	NOR2X1 NOR2X1_1039 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6061), .Y(dp.rf._abc_6362_n9258) );
	NOR2X1 NOR2X1_1040 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9257), .B(dp.rf._abc_6362_n9258), .Y(dp.rf._abc_6362_n9259) );
	NOR2X1 NOR2X1_1041 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9255), .B(dp.rf._abc_6362_n9259), .Y(dp.rf._abc_6362_n9260) );
	NAND2X1 NAND2X1_6273 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9260), .Y(dp.rf._abc_6362_n9261) );
	NAND2X1 NAND2X1_6274 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<7>), .Y(dp.rf._abc_6362_n9262) );
	NAND2X1 NAND2X1_6275 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9262), .Y(dp.rf._abc_6362_n9263) );
	NOR2X1 NOR2X1_1042 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6068), .Y(dp.rf._abc_6362_n9264) );
	NOR2X1 NOR2X1_1043 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9263), .B(dp.rf._abc_6362_n9264), .Y(dp.rf._abc_6362_n9265) );
	NAND2X1 NAND2X1_6276 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<7>), .Y(dp.rf._abc_6362_n9266) );
	NAND2X1 NAND2X1_6277 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9266), .Y(dp.rf._abc_6362_n9267) );
	NOR2X1 NOR2X1_1044 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6073), .Y(dp.rf._abc_6362_n9268) );
	NOR2X1 NOR2X1_1045 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9267), .B(dp.rf._abc_6362_n9268), .Y(dp.rf._abc_6362_n9269) );
	NOR2X1 NOR2X1_1046 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9265), .B(dp.rf._abc_6362_n9269), .Y(dp.rf._abc_6362_n9270) );
	NAND2X1 NAND2X1_6278 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9270), .Y(dp.rf._abc_6362_n9271) );
	NAND2X1 NAND2X1_6279 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9261), .B(dp.rf._abc_6362_n9271), .Y(dp.rf._abc_6362_n9272) );
	NAND2X1 NAND2X1_6280 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9272), .Y(dp.rf._abc_6362_n9273) );
	NAND2X1 NAND2X1_6281 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9273), .Y(dp.rf._abc_6362_n9274) );
	NOR2X1 NOR2X1_1047 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9251), .B(dp.rf._abc_6362_n9274), .Y(dp.rf._abc_6362_n9275) );
	NAND2X1 NAND2X1_6282 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<7>), .Y(dp.rf._abc_6362_n9276) );
	NAND2X1 NAND2X1_6283 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9276), .Y(dp.rf._abc_6362_n9277) );
	NOR2X1 NOR2X1_1048 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6107), .Y(dp.rf._abc_6362_n9278) );
	NOR2X1 NOR2X1_1049 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9277), .B(dp.rf._abc_6362_n9278), .Y(dp.rf._abc_6362_n9279) );
	NAND2X1 NAND2X1_6284 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<7>), .Y(dp.rf._abc_6362_n9280) );
	NAND2X1 NAND2X1_6285 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9280), .Y(dp.rf._abc_6362_n9281) );
	NOR2X1 NOR2X1_1050 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6112), .Y(dp.rf._abc_6362_n9282) );
	NOR2X1 NOR2X1_1051 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9281), .B(dp.rf._abc_6362_n9282), .Y(dp.rf._abc_6362_n9283) );
	OR2X2 OR2X2_92 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9279), .B(dp.rf._abc_6362_n9283), .Y(dp.rf._abc_6362_n9284) );
	NAND2X1 NAND2X1_6286 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9284), .Y(dp.rf._abc_6362_n9285) );
	NAND2X1 NAND2X1_6287 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<7>), .Y(dp.rf._abc_6362_n9286) );
	NAND2X1 NAND2X1_6288 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9286), .Y(dp.rf._abc_6362_n9287) );
	NOR2X1 NOR2X1_1052 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6119), .Y(dp.rf._abc_6362_n9288) );
	NOR2X1 NOR2X1_1053 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9287), .B(dp.rf._abc_6362_n9288), .Y(dp.rf._abc_6362_n9289) );
	NAND2X1 NAND2X1_6289 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<7>), .Y(dp.rf._abc_6362_n9290) );
	NAND2X1 NAND2X1_6290 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9290), .Y(dp.rf._abc_6362_n9291) );
	NOR2X1 NOR2X1_1054 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6124), .Y(dp.rf._abc_6362_n9292) );
	NOR2X1 NOR2X1_1055 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9291), .B(dp.rf._abc_6362_n9292), .Y(dp.rf._abc_6362_n9293) );
	OR2X2 OR2X2_93 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9289), .B(dp.rf._abc_6362_n9293), .Y(dp.rf._abc_6362_n9294) );
	NAND2X1 NAND2X1_6291 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9294), .Y(dp.rf._abc_6362_n9295) );
	AND2X2 AND2X2_406 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9295), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n9296) );
	NAND2X1 NAND2X1_6292 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9285), .B(dp.rf._abc_6362_n9296), .Y(dp.rf._abc_6362_n9297) );
	NAND2X1 NAND2X1_6293 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<7>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9298) );
	NAND2X1 NAND2X1_6294 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<7>), .Y(dp.rf._abc_6362_n9299) );
	AND2X2 AND2X2_407 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9299), .B(instr[17]), .Y(dp.rf._abc_6362_n9300) );
	NAND2X1 NAND2X1_6295 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9298), .B(dp.rf._abc_6362_n9300), .Y(dp.rf._abc_6362_n9301) );
	NAND2X1 NAND2X1_6296 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<7>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9302) );
	NAND2X1 NAND2X1_6297 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<7>), .Y(dp.rf._abc_6362_n9303) );
	AND2X2 AND2X2_408 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9303), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9304) );
	NAND2X1 NAND2X1_6298 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9302), .B(dp.rf._abc_6362_n9304), .Y(dp.rf._abc_6362_n9305) );
	NAND2X1 NAND2X1_6299 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9301), .B(dp.rf._abc_6362_n9305), .Y(dp.rf._abc_6362_n9306) );
	AND2X2 AND2X2_409 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9306), .B(instr[18]), .Y(dp.rf._abc_6362_n9307) );
	NAND2X1 NAND2X1_6300 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<7>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9308) );
	NAND2X1 NAND2X1_6301 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<7>), .Y(dp.rf._abc_6362_n9309) );
	AND2X2 AND2X2_410 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9309), .B(instr[17]), .Y(dp.rf._abc_6362_n9310) );
	NAND2X1 NAND2X1_6302 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9308), .B(dp.rf._abc_6362_n9310), .Y(dp.rf._abc_6362_n9311) );
	NAND2X1 NAND2X1_6303 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<7>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9312) );
	NAND2X1 NAND2X1_6304 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<7>), .Y(dp.rf._abc_6362_n9313) );
	AND2X2 AND2X2_411 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9313), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9314) );
	NAND2X1 NAND2X1_6305 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9312), .B(dp.rf._abc_6362_n9314), .Y(dp.rf._abc_6362_n9315) );
	NAND2X1 NAND2X1_6306 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9311), .B(dp.rf._abc_6362_n9315), .Y(dp.rf._abc_6362_n9316) );
	NAND2X1 NAND2X1_6307 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9316), .Y(dp.rf._abc_6362_n9317) );
	NAND2X1 NAND2X1_6308 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9317), .Y(dp.rf._abc_6362_n9318) );
	NOR2X1 NOR2X1_1056 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9307), .B(dp.rf._abc_6362_n9318), .Y(dp.rf._abc_6362_n9319) );
	NOR2X1 NOR2X1_1057 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9319), .Y(dp.rf._abc_6362_n9320) );
	NAND2X1 NAND2X1_6309 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9297), .B(dp.rf._abc_6362_n9320), .Y(dp.rf._abc_6362_n9321) );
	NAND2X1 NAND2X1_6310 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n9321), .Y(dp.rf._abc_6362_n9322) );
	NOR2X1 NOR2X1_1058 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9275), .B(dp.rf._abc_6362_n9322), .Y(writedata_7__RAW) );
	NAND2X1 NAND2X1_6311 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<8>), .Y(dp.rf._abc_6362_n9324) );
	NAND2X1 NAND2X1_6312 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9324), .Y(dp.rf._abc_6362_n9325) );
	NOR2X1 NOR2X1_1059 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6181), .Y(dp.rf._abc_6362_n9326) );
	NOR2X1 NOR2X1_1060 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9325), .B(dp.rf._abc_6362_n9326), .Y(dp.rf._abc_6362_n9327) );
	NAND2X1 NAND2X1_6313 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<8>), .Y(dp.rf._abc_6362_n9328) );
	NAND2X1 NAND2X1_6314 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9328), .Y(dp.rf._abc_6362_n9329) );
	NOR2X1 NOR2X1_1061 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6186), .Y(dp.rf._abc_6362_n9330) );
	NOR2X1 NOR2X1_1062 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9329), .B(dp.rf._abc_6362_n9330), .Y(dp.rf._abc_6362_n9331) );
	NOR2X1 NOR2X1_1063 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9327), .B(dp.rf._abc_6362_n9331), .Y(dp.rf._abc_6362_n9332) );
	NAND2X1 NAND2X1_6315 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9332), .Y(dp.rf._abc_6362_n9333) );
	NAND2X1 NAND2X1_6316 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<8>), .Y(dp.rf._abc_6362_n9334) );
	NAND2X1 NAND2X1_6317 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9334), .Y(dp.rf._abc_6362_n9335) );
	NOR2X1 NOR2X1_1064 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6193), .Y(dp.rf._abc_6362_n9336) );
	NOR2X1 NOR2X1_1065 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9335), .B(dp.rf._abc_6362_n9336), .Y(dp.rf._abc_6362_n9337) );
	NAND2X1 NAND2X1_6318 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<8>), .Y(dp.rf._abc_6362_n9338) );
	NAND2X1 NAND2X1_6319 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9338), .Y(dp.rf._abc_6362_n9339) );
	NOR2X1 NOR2X1_1066 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6198), .Y(dp.rf._abc_6362_n9340) );
	NOR2X1 NOR2X1_1067 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9339), .B(dp.rf._abc_6362_n9340), .Y(dp.rf._abc_6362_n9341) );
	NOR2X1 NOR2X1_1068 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9337), .B(dp.rf._abc_6362_n9341), .Y(dp.rf._abc_6362_n9342) );
	NAND2X1 NAND2X1_6320 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9342), .Y(dp.rf._abc_6362_n9343) );
	NAND2X1 NAND2X1_6321 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9333), .B(dp.rf._abc_6362_n9343), .Y(dp.rf._abc_6362_n9344) );
	NAND2X1 NAND2X1_6322 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9344), .Y(dp.rf._abc_6362_n9345) );
	NAND2X1 NAND2X1_6323 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<8>), .Y(dp.rf._abc_6362_n9346) );
	NAND2X1 NAND2X1_6324 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<8>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9347) );
	NAND2X1 NAND2X1_6325 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9346), .B(dp.rf._abc_6362_n9347), .Y(dp.rf._abc_6362_n9348) );
	NAND2X1 NAND2X1_6326 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9348), .Y(dp.rf._abc_6362_n9349) );
	NAND2X1 NAND2X1_6327 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<8>), .Y(dp.rf._abc_6362_n9350) );
	NAND2X1 NAND2X1_6328 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<8>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9351) );
	NAND2X1 NAND2X1_6329 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9350), .B(dp.rf._abc_6362_n9351), .Y(dp.rf._abc_6362_n9352) );
	NAND2X1 NAND2X1_6330 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9352), .Y(dp.rf._abc_6362_n9353) );
	AND2X2 AND2X2_412 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9349), .B(dp.rf._abc_6362_n9353), .Y(dp.rf._abc_6362_n9354) );
	NAND2X1 NAND2X1_6331 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9354), .Y(dp.rf._abc_6362_n9355) );
	NAND2X1 NAND2X1_6332 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<8>), .Y(dp.rf._abc_6362_n9356) );
	NAND2X1 NAND2X1_6333 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9356), .Y(dp.rf._abc_6362_n9357) );
	AND2X2 AND2X2_413 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf.rf_2_<8>), .Y(dp.rf._abc_6362_n9358) );
	NOR2X1 NOR2X1_1069 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9357), .B(dp.rf._abc_6362_n9358), .Y(dp.rf._abc_6362_n9359) );
	NAND2X1 NAND2X1_6334 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<8>), .Y(dp.rf._abc_6362_n9360) );
	NAND2X1 NAND2X1_6335 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9360), .Y(dp.rf._abc_6362_n9361) );
	INVX1 INVX1_256 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<8>), .Y(dp.rf._abc_6362_n9362) );
	NOR2X1 NOR2X1_1070 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n9362), .Y(dp.rf._abc_6362_n9363) );
	NOR2X1 NOR2X1_1071 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9361), .B(dp.rf._abc_6362_n9363), .Y(dp.rf._abc_6362_n9364) );
	OR2X2 OR2X2_94 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9359), .B(dp.rf._abc_6362_n9364), .Y(dp.rf._abc_6362_n9365) );
	NAND2X1 NAND2X1_6336 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9365), .Y(dp.rf._abc_6362_n9366) );
	AND2X2 AND2X2_414 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9366), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n9367) );
	NAND2X1 NAND2X1_6337 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9355), .B(dp.rf._abc_6362_n9367), .Y(dp.rf._abc_6362_n9368) );
	NAND2X1 NAND2X1_6338 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9345), .B(dp.rf._abc_6362_n9368), .Y(dp.rf._abc_6362_n9369) );
	NOR2X1 NOR2X1_1072 ( .gnd(gnd), .vdd(vdd), .A(instr[20]), .B(dp.rf._abc_6362_n9369), .Y(dp.rf._abc_6362_n9370) );
	NAND2X1 NAND2X1_6339 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<8>), .Y(dp.rf._abc_6362_n9371) );
	NAND2X1 NAND2X1_6340 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<8>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9372) );
	NAND2X1 NAND2X1_6341 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9371), .B(dp.rf._abc_6362_n9372), .Y(dp.rf._abc_6362_n9373) );
	NAND2X1 NAND2X1_6342 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9373), .Y(dp.rf._abc_6362_n9374) );
	NAND2X1 NAND2X1_6343 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<8>), .Y(dp.rf._abc_6362_n9375) );
	NAND2X1 NAND2X1_6344 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<8>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9376) );
	NAND2X1 NAND2X1_6345 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9375), .B(dp.rf._abc_6362_n9376), .Y(dp.rf._abc_6362_n9377) );
	NAND2X1 NAND2X1_6346 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9377), .Y(dp.rf._abc_6362_n9378) );
	AND2X2 AND2X2_415 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9374), .B(dp.rf._abc_6362_n9378), .Y(dp.rf._abc_6362_n9379) );
	NAND2X1 NAND2X1_6347 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9379), .Y(dp.rf._abc_6362_n9380) );
	NAND2X1 NAND2X1_6348 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<8>), .Y(dp.rf._abc_6362_n9381) );
	NAND2X1 NAND2X1_6349 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<8>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9382) );
	NAND2X1 NAND2X1_6350 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9381), .B(dp.rf._abc_6362_n9382), .Y(dp.rf._abc_6362_n9383) );
	NAND2X1 NAND2X1_6351 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9383), .Y(dp.rf._abc_6362_n9384) );
	NAND2X1 NAND2X1_6352 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<8>), .Y(dp.rf._abc_6362_n9385) );
	NAND2X1 NAND2X1_6353 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<8>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9386) );
	NAND2X1 NAND2X1_6354 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9385), .B(dp.rf._abc_6362_n9386), .Y(dp.rf._abc_6362_n9387) );
	NAND2X1 NAND2X1_6355 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9387), .Y(dp.rf._abc_6362_n9388) );
	AND2X2 AND2X2_416 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9384), .B(dp.rf._abc_6362_n9388), .Y(dp.rf._abc_6362_n9389) );
	NAND2X1 NAND2X1_6356 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9389), .Y(dp.rf._abc_6362_n9390) );
	AND2X2 AND2X2_417 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9390), .B(instr[19]), .Y(dp.rf._abc_6362_n9391) );
	NAND2X1 NAND2X1_6357 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9380), .B(dp.rf._abc_6362_n9391), .Y(dp.rf._abc_6362_n9392) );
	NAND2X1 NAND2X1_6358 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<8>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9393) );
	NAND2X1 NAND2X1_6359 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<8>), .Y(dp.rf._abc_6362_n9394) );
	AND2X2 AND2X2_418 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9394), .B(instr[17]), .Y(dp.rf._abc_6362_n9395) );
	NAND2X1 NAND2X1_6360 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9393), .B(dp.rf._abc_6362_n9395), .Y(dp.rf._abc_6362_n9396) );
	NAND2X1 NAND2X1_6361 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<8>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9397) );
	NAND2X1 NAND2X1_6362 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<8>), .Y(dp.rf._abc_6362_n9398) );
	AND2X2 AND2X2_419 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9398), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9399) );
	NAND2X1 NAND2X1_6363 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9397), .B(dp.rf._abc_6362_n9399), .Y(dp.rf._abc_6362_n9400) );
	NAND2X1 NAND2X1_6364 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9396), .B(dp.rf._abc_6362_n9400), .Y(dp.rf._abc_6362_n9401) );
	AND2X2 AND2X2_420 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9401), .B(instr[18]), .Y(dp.rf._abc_6362_n9402) );
	NAND2X1 NAND2X1_6365 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<8>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9403) );
	NAND2X1 NAND2X1_6366 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<8>), .Y(dp.rf._abc_6362_n9404) );
	AND2X2 AND2X2_421 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9404), .B(instr[17]), .Y(dp.rf._abc_6362_n9405) );
	NAND2X1 NAND2X1_6367 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9403), .B(dp.rf._abc_6362_n9405), .Y(dp.rf._abc_6362_n9406) );
	NAND2X1 NAND2X1_6368 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<8>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9407) );
	NAND2X1 NAND2X1_6369 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<8>), .Y(dp.rf._abc_6362_n9408) );
	AND2X2 AND2X2_422 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9408), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9409) );
	NAND2X1 NAND2X1_6370 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9407), .B(dp.rf._abc_6362_n9409), .Y(dp.rf._abc_6362_n9410) );
	NAND2X1 NAND2X1_6371 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9406), .B(dp.rf._abc_6362_n9410), .Y(dp.rf._abc_6362_n9411) );
	NAND2X1 NAND2X1_6372 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9411), .Y(dp.rf._abc_6362_n9412) );
	NAND2X1 NAND2X1_6373 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n9412), .Y(dp.rf._abc_6362_n9413) );
	NOR2X1 NOR2X1_1073 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9402), .B(dp.rf._abc_6362_n9413), .Y(dp.rf._abc_6362_n9414) );
	NOR2X1 NOR2X1_1074 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9414), .Y(dp.rf._abc_6362_n9415) );
	NAND2X1 NAND2X1_6374 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9392), .B(dp.rf._abc_6362_n9415), .Y(dp.rf._abc_6362_n9416) );
	NAND2X1 NAND2X1_6375 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n9416), .Y(dp.rf._abc_6362_n9417) );
	NOR2X1 NOR2X1_1075 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9370), .B(dp.rf._abc_6362_n9417), .Y(writedata_8__RAW) );
	NAND2X1 NAND2X1_6376 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<9>), .Y(dp.rf._abc_6362_n9419) );
	NAND2X1 NAND2X1_6377 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9419), .Y(dp.rf._abc_6362_n9420) );
	NOR2X1 NOR2X1_1076 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6257), .Y(dp.rf._abc_6362_n9421) );
	NOR2X1 NOR2X1_1077 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9420), .B(dp.rf._abc_6362_n9421), .Y(dp.rf._abc_6362_n9422) );
	NAND2X1 NAND2X1_6378 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<9>), .Y(dp.rf._abc_6362_n9423) );
	NAND2X1 NAND2X1_6379 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9423), .Y(dp.rf._abc_6362_n9424) );
	NOR2X1 NOR2X1_1078 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6262), .Y(dp.rf._abc_6362_n9425) );
	NOR2X1 NOR2X1_1079 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9424), .B(dp.rf._abc_6362_n9425), .Y(dp.rf._abc_6362_n9426) );
	NOR2X1 NOR2X1_1080 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9422), .B(dp.rf._abc_6362_n9426), .Y(dp.rf._abc_6362_n9427) );
	NAND2X1 NAND2X1_6380 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9427), .Y(dp.rf._abc_6362_n9428) );
	NAND2X1 NAND2X1_6381 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<9>), .Y(dp.rf._abc_6362_n9429) );
	NAND2X1 NAND2X1_6382 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9429), .Y(dp.rf._abc_6362_n9430) );
	NOR2X1 NOR2X1_1081 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6269), .Y(dp.rf._abc_6362_n9431) );
	NOR2X1 NOR2X1_1082 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9430), .B(dp.rf._abc_6362_n9431), .Y(dp.rf._abc_6362_n9432) );
	NAND2X1 NAND2X1_6383 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<9>), .Y(dp.rf._abc_6362_n9433) );
	NAND2X1 NAND2X1_6384 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9433), .Y(dp.rf._abc_6362_n9434) );
	NOR2X1 NOR2X1_1083 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6274), .Y(dp.rf._abc_6362_n9435) );
	NOR2X1 NOR2X1_1084 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9434), .B(dp.rf._abc_6362_n9435), .Y(dp.rf._abc_6362_n9436) );
	NOR2X1 NOR2X1_1085 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9432), .B(dp.rf._abc_6362_n9436), .Y(dp.rf._abc_6362_n9437) );
	NAND2X1 NAND2X1_6385 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9437), .Y(dp.rf._abc_6362_n9438) );
	NAND2X1 NAND2X1_6386 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9428), .B(dp.rf._abc_6362_n9438), .Y(dp.rf._abc_6362_n9439) );
	NAND2X1 NAND2X1_6387 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9439), .Y(dp.rf._abc_6362_n9440) );
	NAND2X1 NAND2X1_6388 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<9>), .Y(dp.rf._abc_6362_n9441) );
	NAND2X1 NAND2X1_6389 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9441), .Y(dp.rf._abc_6362_n9442) );
	NOR2X1 NOR2X1_1086 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6283), .Y(dp.rf._abc_6362_n9443) );
	NOR2X1 NOR2X1_1087 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9442), .B(dp.rf._abc_6362_n9443), .Y(dp.rf._abc_6362_n9444) );
	NAND2X1 NAND2X1_6390 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<9>), .Y(dp.rf._abc_6362_n9445) );
	NAND2X1 NAND2X1_6391 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9445), .Y(dp.rf._abc_6362_n9446) );
	NOR2X1 NOR2X1_1088 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6288), .Y(dp.rf._abc_6362_n9447) );
	NOR2X1 NOR2X1_1089 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9446), .B(dp.rf._abc_6362_n9447), .Y(dp.rf._abc_6362_n9448) );
	OR2X2 OR2X2_95 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9444), .B(dp.rf._abc_6362_n9448), .Y(dp.rf._abc_6362_n9449) );
	NAND2X1 NAND2X1_6392 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9449), .Y(dp.rf._abc_6362_n9450) );
	NAND2X1 NAND2X1_6393 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<9>), .Y(dp.rf._abc_6362_n9451) );
	NAND2X1 NAND2X1_6394 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9451), .Y(dp.rf._abc_6362_n9452) );
	NOR2X1 NOR2X1_1090 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6295), .Y(dp.rf._abc_6362_n9453) );
	NOR2X1 NOR2X1_1091 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9452), .B(dp.rf._abc_6362_n9453), .Y(dp.rf._abc_6362_n9454) );
	NAND2X1 NAND2X1_6395 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<9>), .Y(dp.rf._abc_6362_n9455) );
	NAND2X1 NAND2X1_6396 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9455), .Y(dp.rf._abc_6362_n9456) );
	NOR2X1 NOR2X1_1092 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6300), .Y(dp.rf._abc_6362_n9457) );
	NOR2X1 NOR2X1_1093 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9456), .B(dp.rf._abc_6362_n9457), .Y(dp.rf._abc_6362_n9458) );
	OR2X2 OR2X2_96 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9454), .B(dp.rf._abc_6362_n9458), .Y(dp.rf._abc_6362_n9459) );
	NAND2X1 NAND2X1_6397 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9459), .Y(dp.rf._abc_6362_n9460) );
	AND2X2 AND2X2_423 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9460), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n9461) );
	NAND2X1 NAND2X1_6398 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9450), .B(dp.rf._abc_6362_n9461), .Y(dp.rf._abc_6362_n9462) );
	NAND2X1 NAND2X1_6399 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9440), .B(dp.rf._abc_6362_n9462), .Y(dp.rf._abc_6362_n9463) );
	NOR2X1 NOR2X1_1094 ( .gnd(gnd), .vdd(vdd), .A(instr[20]), .B(dp.rf._abc_6362_n9463), .Y(dp.rf._abc_6362_n9464) );
	NAND2X1 NAND2X1_6400 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<9>), .Y(dp.rf._abc_6362_n9465) );
	NAND2X1 NAND2X1_6401 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<9>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9466) );
	NAND2X1 NAND2X1_6402 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9465), .B(dp.rf._abc_6362_n9466), .Y(dp.rf._abc_6362_n9467) );
	NAND2X1 NAND2X1_6403 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9467), .Y(dp.rf._abc_6362_n9468) );
	NAND2X1 NAND2X1_6404 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<9>), .Y(dp.rf._abc_6362_n9469) );
	NAND2X1 NAND2X1_6405 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<9>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9470) );
	NAND2X1 NAND2X1_6406 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9469), .B(dp.rf._abc_6362_n9470), .Y(dp.rf._abc_6362_n9471) );
	NAND2X1 NAND2X1_6407 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9471), .Y(dp.rf._abc_6362_n9472) );
	AND2X2 AND2X2_424 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9468), .B(dp.rf._abc_6362_n9472), .Y(dp.rf._abc_6362_n9473) );
	NAND2X1 NAND2X1_6408 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9473), .Y(dp.rf._abc_6362_n9474) );
	NAND2X1 NAND2X1_6409 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<9>), .Y(dp.rf._abc_6362_n9475) );
	NAND2X1 NAND2X1_6410 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<9>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9476) );
	NAND2X1 NAND2X1_6411 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9475), .B(dp.rf._abc_6362_n9476), .Y(dp.rf._abc_6362_n9477) );
	NAND2X1 NAND2X1_6412 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9477), .Y(dp.rf._abc_6362_n9478) );
	NAND2X1 NAND2X1_6413 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<9>), .Y(dp.rf._abc_6362_n9479) );
	NAND2X1 NAND2X1_6414 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<9>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9480) );
	NAND2X1 NAND2X1_6415 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9479), .B(dp.rf._abc_6362_n9480), .Y(dp.rf._abc_6362_n9481) );
	NAND2X1 NAND2X1_6416 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9481), .Y(dp.rf._abc_6362_n9482) );
	AND2X2 AND2X2_425 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9478), .B(dp.rf._abc_6362_n9482), .Y(dp.rf._abc_6362_n9483) );
	NAND2X1 NAND2X1_6417 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9483), .Y(dp.rf._abc_6362_n9484) );
	AND2X2 AND2X2_426 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9484), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n9485) );
	NAND2X1 NAND2X1_6418 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9474), .B(dp.rf._abc_6362_n9485), .Y(dp.rf._abc_6362_n9486) );
	NAND2X1 NAND2X1_6419 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<9>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9487) );
	NAND2X1 NAND2X1_6420 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<9>), .Y(dp.rf._abc_6362_n9488) );
	AND2X2 AND2X2_427 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9488), .B(instr[17]), .Y(dp.rf._abc_6362_n9489) );
	NAND2X1 NAND2X1_6421 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9487), .B(dp.rf._abc_6362_n9489), .Y(dp.rf._abc_6362_n9490) );
	NAND2X1 NAND2X1_6422 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<9>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9491) );
	NAND2X1 NAND2X1_6423 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<9>), .Y(dp.rf._abc_6362_n9492) );
	AND2X2 AND2X2_428 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9492), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9493) );
	NAND2X1 NAND2X1_6424 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9491), .B(dp.rf._abc_6362_n9493), .Y(dp.rf._abc_6362_n9494) );
	NAND2X1 NAND2X1_6425 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9490), .B(dp.rf._abc_6362_n9494), .Y(dp.rf._abc_6362_n9495) );
	AND2X2 AND2X2_429 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9495), .B(instr[18]), .Y(dp.rf._abc_6362_n9496) );
	NAND2X1 NAND2X1_6426 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<9>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9497) );
	NAND2X1 NAND2X1_6427 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<9>), .Y(dp.rf._abc_6362_n9498) );
	AND2X2 AND2X2_430 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9498), .B(instr[17]), .Y(dp.rf._abc_6362_n9499) );
	NAND2X1 NAND2X1_6428 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9497), .B(dp.rf._abc_6362_n9499), .Y(dp.rf._abc_6362_n9500) );
	NAND2X1 NAND2X1_6429 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<9>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9501) );
	NAND2X1 NAND2X1_6430 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<9>), .Y(dp.rf._abc_6362_n9502) );
	AND2X2 AND2X2_431 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9502), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9503) );
	NAND2X1 NAND2X1_6431 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9501), .B(dp.rf._abc_6362_n9503), .Y(dp.rf._abc_6362_n9504) );
	NAND2X1 NAND2X1_6432 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9500), .B(dp.rf._abc_6362_n9504), .Y(dp.rf._abc_6362_n9505) );
	NAND2X1 NAND2X1_6433 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9505), .Y(dp.rf._abc_6362_n9506) );
	NAND2X1 NAND2X1_6434 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9506), .Y(dp.rf._abc_6362_n9507) );
	NOR2X1 NOR2X1_1095 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9496), .B(dp.rf._abc_6362_n9507), .Y(dp.rf._abc_6362_n9508) );
	NOR2X1 NOR2X1_1096 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9508), .Y(dp.rf._abc_6362_n9509) );
	NAND2X1 NAND2X1_6435 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9486), .B(dp.rf._abc_6362_n9509), .Y(dp.rf._abc_6362_n9510) );
	NAND2X1 NAND2X1_6436 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n9510), .Y(dp.rf._abc_6362_n9511) );
	NOR2X1 NOR2X1_1097 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9464), .B(dp.rf._abc_6362_n9511), .Y(writedata_9__RAW) );
	NAND2X1 NAND2X1_6437 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<10>), .Y(dp.rf._abc_6362_n9513) );
	NAND2X1 NAND2X1_6438 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<10>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9514) );
	NAND2X1 NAND2X1_6439 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9513), .B(dp.rf._abc_6362_n9514), .Y(dp.rf._abc_6362_n9515) );
	NAND2X1 NAND2X1_6440 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9515), .Y(dp.rf._abc_6362_n9516) );
	NAND2X1 NAND2X1_6441 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<10>), .Y(dp.rf._abc_6362_n9517) );
	NAND2X1 NAND2X1_6442 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<10>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9518) );
	NAND2X1 NAND2X1_6443 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9517), .B(dp.rf._abc_6362_n9518), .Y(dp.rf._abc_6362_n9519) );
	NAND2X1 NAND2X1_6444 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9519), .Y(dp.rf._abc_6362_n9520) );
	NAND2X1 NAND2X1_6445 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9516), .B(dp.rf._abc_6362_n9520), .Y(dp.rf._abc_6362_n9521) );
	NOR2X1 NOR2X1_1098 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9521), .Y(dp.rf._abc_6362_n9522) );
	NAND2X1 NAND2X1_6446 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<10>), .Y(dp.rf._abc_6362_n9523) );
	NAND2X1 NAND2X1_6447 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<10>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9524) );
	NAND2X1 NAND2X1_6448 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9523), .B(dp.rf._abc_6362_n9524), .Y(dp.rf._abc_6362_n9525) );
	NAND2X1 NAND2X1_6449 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9525), .Y(dp.rf._abc_6362_n9526) );
	NAND2X1 NAND2X1_6450 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<10>), .Y(dp.rf._abc_6362_n9527) );
	NAND2X1 NAND2X1_6451 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<10>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9528) );
	NAND2X1 NAND2X1_6452 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9527), .B(dp.rf._abc_6362_n9528), .Y(dp.rf._abc_6362_n9529) );
	NAND2X1 NAND2X1_6453 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9529), .Y(dp.rf._abc_6362_n9530) );
	AND2X2 AND2X2_432 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9526), .B(dp.rf._abc_6362_n9530), .Y(dp.rf._abc_6362_n9531) );
	NAND2X1 NAND2X1_6454 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9531), .Y(dp.rf._abc_6362_n9532) );
	NAND2X1 NAND2X1_6455 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n9532), .Y(dp.rf._abc_6362_n9533) );
	NOR2X1 NOR2X1_1099 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9522), .B(dp.rf._abc_6362_n9533), .Y(dp.rf._abc_6362_n9534) );
	NAND2X1 NAND2X1_6456 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<10>), .Y(dp.rf._abc_6362_n9535) );
	NAND2X1 NAND2X1_6457 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9535), .Y(dp.rf._abc_6362_n9536) );
	NOR2X1 NOR2X1_1100 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6359), .Y(dp.rf._abc_6362_n9537) );
	NOR2X1 NOR2X1_1101 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9536), .B(dp.rf._abc_6362_n9537), .Y(dp.rf._abc_6362_n9538) );
	NAND2X1 NAND2X1_6458 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<10>), .Y(dp.rf._abc_6362_n9539) );
	NAND2X1 NAND2X1_6459 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9539), .Y(dp.rf._abc_6362_n9540) );
	NOR2X1 NOR2X1_1102 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6364), .Y(dp.rf._abc_6362_n9541) );
	NOR2X1 NOR2X1_1103 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9540), .B(dp.rf._abc_6362_n9541), .Y(dp.rf._abc_6362_n9542) );
	NOR2X1 NOR2X1_1104 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9538), .B(dp.rf._abc_6362_n9542), .Y(dp.rf._abc_6362_n9543) );
	NAND2X1 NAND2X1_6460 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9543), .Y(dp.rf._abc_6362_n9544) );
	NAND2X1 NAND2X1_6461 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<10>), .Y(dp.rf._abc_6362_n9545) );
	NAND2X1 NAND2X1_6462 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9545), .Y(dp.rf._abc_6362_n9546) );
	NOR2X1 NOR2X1_1105 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6371), .Y(dp.rf._abc_6362_n9547) );
	NOR2X1 NOR2X1_1106 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9546), .B(dp.rf._abc_6362_n9547), .Y(dp.rf._abc_6362_n9548) );
	NAND2X1 NAND2X1_6463 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<10>), .Y(dp.rf._abc_6362_n9549) );
	NAND2X1 NAND2X1_6464 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9549), .Y(dp.rf._abc_6362_n9550) );
	NOR2X1 NOR2X1_1107 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6376), .Y(dp.rf._abc_6362_n9551) );
	NOR2X1 NOR2X1_1108 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9550), .B(dp.rf._abc_6362_n9551), .Y(dp.rf._abc_6362_n9552) );
	NOR2X1 NOR2X1_1109 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9548), .B(dp.rf._abc_6362_n9552), .Y(dp.rf._abc_6362_n9553) );
	NAND2X1 NAND2X1_6465 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9553), .Y(dp.rf._abc_6362_n9554) );
	NAND2X1 NAND2X1_6466 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9544), .B(dp.rf._abc_6362_n9554), .Y(dp.rf._abc_6362_n9555) );
	NAND2X1 NAND2X1_6467 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9555), .Y(dp.rf._abc_6362_n9556) );
	NAND2X1 NAND2X1_6468 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9556), .Y(dp.rf._abc_6362_n9557) );
	NOR2X1 NOR2X1_1110 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9534), .B(dp.rf._abc_6362_n9557), .Y(dp.rf._abc_6362_n9558) );
	NAND2X1 NAND2X1_6469 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<10>), .Y(dp.rf._abc_6362_n9559) );
	NAND2X1 NAND2X1_6470 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9559), .Y(dp.rf._abc_6362_n9560) );
	NOR2X1 NOR2X1_1111 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6410), .Y(dp.rf._abc_6362_n9561) );
	NOR2X1 NOR2X1_1112 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9560), .B(dp.rf._abc_6362_n9561), .Y(dp.rf._abc_6362_n9562) );
	NAND2X1 NAND2X1_6471 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<10>), .Y(dp.rf._abc_6362_n9563) );
	NAND2X1 NAND2X1_6472 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9563), .Y(dp.rf._abc_6362_n9564) );
	NOR2X1 NOR2X1_1113 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6415), .Y(dp.rf._abc_6362_n9565) );
	NOR2X1 NOR2X1_1114 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9564), .B(dp.rf._abc_6362_n9565), .Y(dp.rf._abc_6362_n9566) );
	OR2X2 OR2X2_97 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9562), .B(dp.rf._abc_6362_n9566), .Y(dp.rf._abc_6362_n9567) );
	NAND2X1 NAND2X1_6473 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9567), .Y(dp.rf._abc_6362_n9568) );
	NAND2X1 NAND2X1_6474 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<10>), .Y(dp.rf._abc_6362_n9569) );
	NAND2X1 NAND2X1_6475 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9569), .Y(dp.rf._abc_6362_n9570) );
	NOR2X1 NOR2X1_1115 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6422), .Y(dp.rf._abc_6362_n9571) );
	NOR2X1 NOR2X1_1116 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9570), .B(dp.rf._abc_6362_n9571), .Y(dp.rf._abc_6362_n9572) );
	NAND2X1 NAND2X1_6476 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<10>), .Y(dp.rf._abc_6362_n9573) );
	NAND2X1 NAND2X1_6477 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9573), .Y(dp.rf._abc_6362_n9574) );
	NOR2X1 NOR2X1_1117 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6427), .Y(dp.rf._abc_6362_n9575) );
	NOR2X1 NOR2X1_1118 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9574), .B(dp.rf._abc_6362_n9575), .Y(dp.rf._abc_6362_n9576) );
	OR2X2 OR2X2_98 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9572), .B(dp.rf._abc_6362_n9576), .Y(dp.rf._abc_6362_n9577) );
	NAND2X1 NAND2X1_6478 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9577), .Y(dp.rf._abc_6362_n9578) );
	AND2X2 AND2X2_433 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9578), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n9579) );
	NAND2X1 NAND2X1_6479 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9568), .B(dp.rf._abc_6362_n9579), .Y(dp.rf._abc_6362_n9580) );
	NAND2X1 NAND2X1_6480 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<10>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9581) );
	NAND2X1 NAND2X1_6481 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<10>), .Y(dp.rf._abc_6362_n9582) );
	AND2X2 AND2X2_434 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9582), .B(instr[17]), .Y(dp.rf._abc_6362_n9583) );
	NAND2X1 NAND2X1_6482 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9581), .B(dp.rf._abc_6362_n9583), .Y(dp.rf._abc_6362_n9584) );
	NAND2X1 NAND2X1_6483 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<10>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9585) );
	NAND2X1 NAND2X1_6484 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<10>), .Y(dp.rf._abc_6362_n9586) );
	AND2X2 AND2X2_435 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9586), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9587) );
	NAND2X1 NAND2X1_6485 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9585), .B(dp.rf._abc_6362_n9587), .Y(dp.rf._abc_6362_n9588) );
	NAND2X1 NAND2X1_6486 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9584), .B(dp.rf._abc_6362_n9588), .Y(dp.rf._abc_6362_n9589) );
	AND2X2 AND2X2_436 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9589), .B(instr[18]), .Y(dp.rf._abc_6362_n9590) );
	NAND2X1 NAND2X1_6487 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<10>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9591) );
	NAND2X1 NAND2X1_6488 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<10>), .Y(dp.rf._abc_6362_n9592) );
	AND2X2 AND2X2_437 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9592), .B(instr[17]), .Y(dp.rf._abc_6362_n9593) );
	NAND2X1 NAND2X1_6489 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9591), .B(dp.rf._abc_6362_n9593), .Y(dp.rf._abc_6362_n9594) );
	NAND2X1 NAND2X1_6490 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<10>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9595) );
	NAND2X1 NAND2X1_6491 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<10>), .Y(dp.rf._abc_6362_n9596) );
	AND2X2 AND2X2_438 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9596), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9597) );
	NAND2X1 NAND2X1_6492 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9595), .B(dp.rf._abc_6362_n9597), .Y(dp.rf._abc_6362_n9598) );
	NAND2X1 NAND2X1_6493 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9594), .B(dp.rf._abc_6362_n9598), .Y(dp.rf._abc_6362_n9599) );
	NAND2X1 NAND2X1_6494 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9599), .Y(dp.rf._abc_6362_n9600) );
	NAND2X1 NAND2X1_6495 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9600), .Y(dp.rf._abc_6362_n9601) );
	NOR2X1 NOR2X1_1119 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9590), .B(dp.rf._abc_6362_n9601), .Y(dp.rf._abc_6362_n9602) );
	NOR2X1 NOR2X1_1120 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9602), .Y(dp.rf._abc_6362_n9603) );
	NAND2X1 NAND2X1_6496 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9580), .B(dp.rf._abc_6362_n9603), .Y(dp.rf._abc_6362_n9604) );
	NAND2X1 NAND2X1_6497 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n9604), .Y(dp.rf._abc_6362_n9605) );
	NOR2X1 NOR2X1_1121 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9558), .B(dp.rf._abc_6362_n9605), .Y(writedata_10__RAW) );
	NAND2X1 NAND2X1_6498 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<11>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9607) );
	NOR2X1 NOR2X1_1122 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6488), .Y(dp.rf._abc_6362_n9608) );
	NOR2X1 NOR2X1_1123 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9608), .Y(dp.rf._abc_6362_n9609) );
	NAND2X1 NAND2X1_6499 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9607), .B(dp.rf._abc_6362_n9609), .Y(dp.rf._abc_6362_n9610) );
	NAND2X1 NAND2X1_6500 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<11>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9611) );
	NOR2X1 NOR2X1_1124 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6493), .Y(dp.rf._abc_6362_n9612) );
	NOR2X1 NOR2X1_1125 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9612), .Y(dp.rf._abc_6362_n9613) );
	NAND2X1 NAND2X1_6501 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9611), .B(dp.rf._abc_6362_n9613), .Y(dp.rf._abc_6362_n9614) );
	NAND2X1 NAND2X1_6502 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9610), .B(dp.rf._abc_6362_n9614), .Y(dp.rf._abc_6362_n9615) );
	NOR2X1 NOR2X1_1126 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9615), .Y(dp.rf._abc_6362_n9616) );
	NAND2X1 NAND2X1_6503 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<11>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9617) );
	NOR2X1 NOR2X1_1127 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6500), .Y(dp.rf._abc_6362_n9618) );
	NOR2X1 NOR2X1_1128 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9618), .Y(dp.rf._abc_6362_n9619) );
	NAND2X1 NAND2X1_6504 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9617), .B(dp.rf._abc_6362_n9619), .Y(dp.rf._abc_6362_n9620) );
	NAND2X1 NAND2X1_6505 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<11>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9621) );
	NOR2X1 NOR2X1_1129 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6505), .Y(dp.rf._abc_6362_n9622) );
	NOR2X1 NOR2X1_1130 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9622), .Y(dp.rf._abc_6362_n9623) );
	NAND2X1 NAND2X1_6506 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9621), .B(dp.rf._abc_6362_n9623), .Y(dp.rf._abc_6362_n9624) );
	NAND2X1 NAND2X1_6507 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9620), .B(dp.rf._abc_6362_n9624), .Y(dp.rf._abc_6362_n9625) );
	NOR2X1 NOR2X1_1131 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9625), .Y(dp.rf._abc_6362_n9626) );
	NOR2X1 NOR2X1_1132 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9616), .B(dp.rf._abc_6362_n9626), .Y(dp.rf._abc_6362_n9627) );
	NOR2X1 NOR2X1_1133 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9627), .Y(dp.rf._abc_6362_n9628) );
	NAND2X1 NAND2X1_6508 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<11>), .Y(dp.rf._abc_6362_n9629) );
	NAND2X1 NAND2X1_6509 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9629), .Y(dp.rf._abc_6362_n9630) );
	NOR2X1 NOR2X1_1134 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6474), .Y(dp.rf._abc_6362_n9631) );
	NOR2X1 NOR2X1_1135 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9630), .B(dp.rf._abc_6362_n9631), .Y(dp.rf._abc_6362_n9632) );
	NAND2X1 NAND2X1_6510 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<11>), .Y(dp.rf._abc_6362_n9633) );
	NAND2X1 NAND2X1_6511 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9633), .Y(dp.rf._abc_6362_n9634) );
	NOR2X1 NOR2X1_1136 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6479), .Y(dp.rf._abc_6362_n9635) );
	NOR2X1 NOR2X1_1137 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9634), .B(dp.rf._abc_6362_n9635), .Y(dp.rf._abc_6362_n9636) );
	OR2X2 OR2X2_99 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9632), .B(dp.rf._abc_6362_n9636), .Y(dp.rf._abc_6362_n9637) );
	NAND2X1 NAND2X1_6512 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9637), .Y(dp.rf._abc_6362_n9638) );
	NAND2X1 NAND2X1_6513 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<11>), .Y(dp.rf._abc_6362_n9639) );
	NAND2X1 NAND2X1_6514 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9639), .Y(dp.rf._abc_6362_n9640) );
	NOR2X1 NOR2X1_1138 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6462), .Y(dp.rf._abc_6362_n9641) );
	NOR2X1 NOR2X1_1139 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9640), .B(dp.rf._abc_6362_n9641), .Y(dp.rf._abc_6362_n9642) );
	NAND2X1 NAND2X1_6515 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<11>), .Y(dp.rf._abc_6362_n9643) );
	NAND2X1 NAND2X1_6516 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9643), .Y(dp.rf._abc_6362_n9644) );
	NOR2X1 NOR2X1_1140 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6467), .Y(dp.rf._abc_6362_n9645) );
	NOR2X1 NOR2X1_1141 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9644), .B(dp.rf._abc_6362_n9645), .Y(dp.rf._abc_6362_n9646) );
	OR2X2 OR2X2_100 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9642), .B(dp.rf._abc_6362_n9646), .Y(dp.rf._abc_6362_n9647) );
	NAND2X1 NAND2X1_6517 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9647), .Y(dp.rf._abc_6362_n9648) );
	AND2X2 AND2X2_439 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9648), .B(instr[19]), .Y(dp.rf._abc_6362_n9649) );
	NAND2X1 NAND2X1_6518 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9638), .B(dp.rf._abc_6362_n9649), .Y(dp.rf._abc_6362_n9650) );
	NAND2X1 NAND2X1_6519 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9650), .Y(dp.rf._abc_6362_n9651) );
	NOR2X1 NOR2X1_1142 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9628), .B(dp.rf._abc_6362_n9651), .Y(dp.rf._abc_6362_n9652) );
	NAND2X1 NAND2X1_6520 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<11>), .Y(dp.rf._abc_6362_n9653) );
	NAND2X1 NAND2X1_6521 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9653), .Y(dp.rf._abc_6362_n9654) );
	NOR2X1 NOR2X1_1143 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6516), .Y(dp.rf._abc_6362_n9655) );
	NOR2X1 NOR2X1_1144 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9654), .B(dp.rf._abc_6362_n9655), .Y(dp.rf._abc_6362_n9656) );
	NAND2X1 NAND2X1_6522 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<11>), .Y(dp.rf._abc_6362_n9657) );
	NAND2X1 NAND2X1_6523 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9657), .Y(dp.rf._abc_6362_n9658) );
	NOR2X1 NOR2X1_1145 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6521), .Y(dp.rf._abc_6362_n9659) );
	NOR2X1 NOR2X1_1146 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9658), .B(dp.rf._abc_6362_n9659), .Y(dp.rf._abc_6362_n9660) );
	OR2X2 OR2X2_101 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9656), .B(dp.rf._abc_6362_n9660), .Y(dp.rf._abc_6362_n9661) );
	NAND2X1 NAND2X1_6524 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9661), .Y(dp.rf._abc_6362_n9662) );
	NAND2X1 NAND2X1_6525 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<11>), .Y(dp.rf._abc_6362_n9663) );
	NAND2X1 NAND2X1_6526 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9663), .Y(dp.rf._abc_6362_n9664) );
	NOR2X1 NOR2X1_1147 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6528), .Y(dp.rf._abc_6362_n9665) );
	NOR2X1 NOR2X1_1148 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9664), .B(dp.rf._abc_6362_n9665), .Y(dp.rf._abc_6362_n9666) );
	NAND2X1 NAND2X1_6527 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<11>), .Y(dp.rf._abc_6362_n9667) );
	NAND2X1 NAND2X1_6528 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9667), .Y(dp.rf._abc_6362_n9668) );
	NOR2X1 NOR2X1_1149 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6533), .Y(dp.rf._abc_6362_n9669) );
	NOR2X1 NOR2X1_1150 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9668), .B(dp.rf._abc_6362_n9669), .Y(dp.rf._abc_6362_n9670) );
	OR2X2 OR2X2_102 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9666), .B(dp.rf._abc_6362_n9670), .Y(dp.rf._abc_6362_n9671) );
	NAND2X1 NAND2X1_6529 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9671), .Y(dp.rf._abc_6362_n9672) );
	AND2X2 AND2X2_440 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9672), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n9673) );
	NAND2X1 NAND2X1_6530 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9662), .B(dp.rf._abc_6362_n9673), .Y(dp.rf._abc_6362_n9674) );
	NAND2X1 NAND2X1_6531 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<11>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9675) );
	NAND2X1 NAND2X1_6532 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<11>), .Y(dp.rf._abc_6362_n9676) );
	AND2X2 AND2X2_441 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9676), .B(instr[17]), .Y(dp.rf._abc_6362_n9677) );
	NAND2X1 NAND2X1_6533 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9675), .B(dp.rf._abc_6362_n9677), .Y(dp.rf._abc_6362_n9678) );
	NAND2X1 NAND2X1_6534 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<11>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9679) );
	NAND2X1 NAND2X1_6535 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<11>), .Y(dp.rf._abc_6362_n9680) );
	AND2X2 AND2X2_442 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9680), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9681) );
	NAND2X1 NAND2X1_6536 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9679), .B(dp.rf._abc_6362_n9681), .Y(dp.rf._abc_6362_n9682) );
	NAND2X1 NAND2X1_6537 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9678), .B(dp.rf._abc_6362_n9682), .Y(dp.rf._abc_6362_n9683) );
	AND2X2 AND2X2_443 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9683), .B(instr[18]), .Y(dp.rf._abc_6362_n9684) );
	NAND2X1 NAND2X1_6538 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<11>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9685) );
	NAND2X1 NAND2X1_6539 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<11>), .Y(dp.rf._abc_6362_n9686) );
	AND2X2 AND2X2_444 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9686), .B(instr[17]), .Y(dp.rf._abc_6362_n9687) );
	NAND2X1 NAND2X1_6540 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9685), .B(dp.rf._abc_6362_n9687), .Y(dp.rf._abc_6362_n9688) );
	NAND2X1 NAND2X1_6541 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<11>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9689) );
	NAND2X1 NAND2X1_6542 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<11>), .Y(dp.rf._abc_6362_n9690) );
	AND2X2 AND2X2_445 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9690), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9691) );
	NAND2X1 NAND2X1_6543 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9689), .B(dp.rf._abc_6362_n9691), .Y(dp.rf._abc_6362_n9692) );
	NAND2X1 NAND2X1_6544 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9688), .B(dp.rf._abc_6362_n9692), .Y(dp.rf._abc_6362_n9693) );
	NAND2X1 NAND2X1_6545 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9693), .Y(dp.rf._abc_6362_n9694) );
	NAND2X1 NAND2X1_6546 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9694), .Y(dp.rf._abc_6362_n9695) );
	NOR2X1 NOR2X1_1151 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9684), .B(dp.rf._abc_6362_n9695), .Y(dp.rf._abc_6362_n9696) );
	NOR2X1 NOR2X1_1152 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9696), .Y(dp.rf._abc_6362_n9697) );
	NAND2X1 NAND2X1_6547 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9674), .B(dp.rf._abc_6362_n9697), .Y(dp.rf._abc_6362_n9698) );
	NAND2X1 NAND2X1_6548 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n9698), .Y(dp.rf._abc_6362_n9699) );
	NOR2X1 NOR2X1_1153 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9652), .B(dp.rf._abc_6362_n9699), .Y(writedata_11__RAW) );
	NAND2X1 NAND2X1_6549 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<12>), .Y(dp.rf._abc_6362_n9701) );
	NAND2X1 NAND2X1_6550 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9701), .Y(dp.rf._abc_6362_n9702) );
	NOR2X1 NOR2X1_1154 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6606), .Y(dp.rf._abc_6362_n9703) );
	NOR2X1 NOR2X1_1155 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9702), .B(dp.rf._abc_6362_n9703), .Y(dp.rf._abc_6362_n9704) );
	NAND2X1 NAND2X1_6551 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<12>), .Y(dp.rf._abc_6362_n9705) );
	NAND2X1 NAND2X1_6552 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9705), .Y(dp.rf._abc_6362_n9706) );
	NOR2X1 NOR2X1_1156 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6611), .Y(dp.rf._abc_6362_n9707) );
	NOR2X1 NOR2X1_1157 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9706), .B(dp.rf._abc_6362_n9707), .Y(dp.rf._abc_6362_n9708) );
	NOR2X1 NOR2X1_1158 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9704), .B(dp.rf._abc_6362_n9708), .Y(dp.rf._abc_6362_n9709) );
	NAND2X1 NAND2X1_6553 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9709), .Y(dp.rf._abc_6362_n9710) );
	NAND2X1 NAND2X1_6554 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<12>), .Y(dp.rf._abc_6362_n9711) );
	NAND2X1 NAND2X1_6555 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9711), .Y(dp.rf._abc_6362_n9712) );
	NOR2X1 NOR2X1_1159 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6594), .Y(dp.rf._abc_6362_n9713) );
	NOR2X1 NOR2X1_1160 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9712), .B(dp.rf._abc_6362_n9713), .Y(dp.rf._abc_6362_n9714) );
	NAND2X1 NAND2X1_6556 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<12>), .Y(dp.rf._abc_6362_n9715) );
	NAND2X1 NAND2X1_6557 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9715), .Y(dp.rf._abc_6362_n9716) );
	NOR2X1 NOR2X1_1161 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6599), .Y(dp.rf._abc_6362_n9717) );
	NOR2X1 NOR2X1_1162 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9716), .B(dp.rf._abc_6362_n9717), .Y(dp.rf._abc_6362_n9718) );
	NOR2X1 NOR2X1_1163 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9714), .B(dp.rf._abc_6362_n9718), .Y(dp.rf._abc_6362_n9719) );
	NAND2X1 NAND2X1_6558 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9719), .Y(dp.rf._abc_6362_n9720) );
	NAND2X1 NAND2X1_6559 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9710), .B(dp.rf._abc_6362_n9720), .Y(dp.rf._abc_6362_n9721) );
	NAND2X1 NAND2X1_6560 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9721), .Y(dp.rf._abc_6362_n9722) );
	NAND2X1 NAND2X1_6561 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9722), .Y(dp.rf._abc_6362_n9723) );
	NAND2X1 NAND2X1_6562 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9724) );
	NOR2X1 NOR2X1_1164 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6567), .Y(dp.rf._abc_6362_n9725) );
	NOR2X1 NOR2X1_1165 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9725), .Y(dp.rf._abc_6362_n9726) );
	NAND2X1 NAND2X1_6563 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9724), .B(dp.rf._abc_6362_n9726), .Y(dp.rf._abc_6362_n9727) );
	NAND2X1 NAND2X1_6564 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9728) );
	NOR2X1 NOR2X1_1166 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6572), .Y(dp.rf._abc_6362_n9729) );
	NOR2X1 NOR2X1_1167 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9729), .Y(dp.rf._abc_6362_n9730) );
	NAND2X1 NAND2X1_6565 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9728), .B(dp.rf._abc_6362_n9730), .Y(dp.rf._abc_6362_n9731) );
	NAND2X1 NAND2X1_6566 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9727), .B(dp.rf._abc_6362_n9731), .Y(dp.rf._abc_6362_n9732) );
	NOR2X1 NOR2X1_1168 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9732), .Y(dp.rf._abc_6362_n9733) );
	NAND2X1 NAND2X1_6567 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9734) );
	NOR2X1 NOR2X1_1169 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6579), .Y(dp.rf._abc_6362_n9735) );
	NOR2X1 NOR2X1_1170 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9735), .Y(dp.rf._abc_6362_n9736) );
	NAND2X1 NAND2X1_6568 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9734), .B(dp.rf._abc_6362_n9736), .Y(dp.rf._abc_6362_n9737) );
	NAND2X1 NAND2X1_6569 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9738) );
	NOR2X1 NOR2X1_1171 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6584), .Y(dp.rf._abc_6362_n9739) );
	NOR2X1 NOR2X1_1172 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9739), .Y(dp.rf._abc_6362_n9740) );
	NAND2X1 NAND2X1_6570 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9738), .B(dp.rf._abc_6362_n9740), .Y(dp.rf._abc_6362_n9741) );
	NAND2X1 NAND2X1_6571 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9737), .B(dp.rf._abc_6362_n9741), .Y(dp.rf._abc_6362_n9742) );
	NOR2X1 NOR2X1_1173 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9742), .Y(dp.rf._abc_6362_n9743) );
	NOR2X1 NOR2X1_1174 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9733), .B(dp.rf._abc_6362_n9743), .Y(dp.rf._abc_6362_n9744) );
	NOR2X1 NOR2X1_1175 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9744), .Y(dp.rf._abc_6362_n9745) );
	NOR2X1 NOR2X1_1176 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9723), .B(dp.rf._abc_6362_n9745), .Y(dp.rf._abc_6362_n9746) );
	NAND2X1 NAND2X1_6572 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<12>), .Y(dp.rf._abc_6362_n9747) );
	NAND2X1 NAND2X1_6573 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9748) );
	NAND2X1 NAND2X1_6574 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9747), .B(dp.rf._abc_6362_n9748), .Y(dp.rf._abc_6362_n9749) );
	NAND2X1 NAND2X1_6575 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9749), .Y(dp.rf._abc_6362_n9750) );
	NAND2X1 NAND2X1_6576 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<12>), .Y(dp.rf._abc_6362_n9751) );
	NAND2X1 NAND2X1_6577 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9752) );
	NAND2X1 NAND2X1_6578 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9751), .B(dp.rf._abc_6362_n9752), .Y(dp.rf._abc_6362_n9753) );
	NAND2X1 NAND2X1_6579 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9753), .Y(dp.rf._abc_6362_n9754) );
	AND2X2 AND2X2_446 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9750), .B(dp.rf._abc_6362_n9754), .Y(dp.rf._abc_6362_n9755) );
	NAND2X1 NAND2X1_6580 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9755), .Y(dp.rf._abc_6362_n9756) );
	NAND2X1 NAND2X1_6581 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<12>), .Y(dp.rf._abc_6362_n9757) );
	NAND2X1 NAND2X1_6582 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9758) );
	NAND2X1 NAND2X1_6583 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9757), .B(dp.rf._abc_6362_n9758), .Y(dp.rf._abc_6362_n9759) );
	NAND2X1 NAND2X1_6584 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9759), .Y(dp.rf._abc_6362_n9760) );
	NAND2X1 NAND2X1_6585 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<12>), .Y(dp.rf._abc_6362_n9761) );
	NAND2X1 NAND2X1_6586 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9762) );
	NAND2X1 NAND2X1_6587 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9761), .B(dp.rf._abc_6362_n9762), .Y(dp.rf._abc_6362_n9763) );
	NAND2X1 NAND2X1_6588 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9763), .Y(dp.rf._abc_6362_n9764) );
	AND2X2 AND2X2_447 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9760), .B(dp.rf._abc_6362_n9764), .Y(dp.rf._abc_6362_n9765) );
	NAND2X1 NAND2X1_6589 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9765), .Y(dp.rf._abc_6362_n9766) );
	AND2X2 AND2X2_448 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9766), .B(instr[19]), .Y(dp.rf._abc_6362_n9767) );
	NAND2X1 NAND2X1_6590 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9756), .B(dp.rf._abc_6362_n9767), .Y(dp.rf._abc_6362_n9768) );
	NAND2X1 NAND2X1_6591 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9769) );
	NAND2X1 NAND2X1_6592 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<12>), .Y(dp.rf._abc_6362_n9770) );
	AND2X2 AND2X2_449 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9770), .B(instr[17]), .Y(dp.rf._abc_6362_n9771) );
	NAND2X1 NAND2X1_6593 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9769), .B(dp.rf._abc_6362_n9771), .Y(dp.rf._abc_6362_n9772) );
	NAND2X1 NAND2X1_6594 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9773) );
	NAND2X1 NAND2X1_6595 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<12>), .Y(dp.rf._abc_6362_n9774) );
	AND2X2 AND2X2_450 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9774), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9775) );
	NAND2X1 NAND2X1_6596 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9773), .B(dp.rf._abc_6362_n9775), .Y(dp.rf._abc_6362_n9776) );
	NAND2X1 NAND2X1_6597 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9772), .B(dp.rf._abc_6362_n9776), .Y(dp.rf._abc_6362_n9777) );
	AND2X2 AND2X2_451 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9777), .B(instr[18]), .Y(dp.rf._abc_6362_n9778) );
	NAND2X1 NAND2X1_6598 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9779) );
	NAND2X1 NAND2X1_6599 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<12>), .Y(dp.rf._abc_6362_n9780) );
	AND2X2 AND2X2_452 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9780), .B(instr[17]), .Y(dp.rf._abc_6362_n9781) );
	NAND2X1 NAND2X1_6600 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9779), .B(dp.rf._abc_6362_n9781), .Y(dp.rf._abc_6362_n9782) );
	NAND2X1 NAND2X1_6601 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<12>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9783) );
	NAND2X1 NAND2X1_6602 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<12>), .Y(dp.rf._abc_6362_n9784) );
	AND2X2 AND2X2_453 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9784), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9785) );
	NAND2X1 NAND2X1_6603 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9783), .B(dp.rf._abc_6362_n9785), .Y(dp.rf._abc_6362_n9786) );
	NAND2X1 NAND2X1_6604 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9782), .B(dp.rf._abc_6362_n9786), .Y(dp.rf._abc_6362_n9787) );
	NAND2X1 NAND2X1_6605 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9787), .Y(dp.rf._abc_6362_n9788) );
	NAND2X1 NAND2X1_6606 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n9788), .Y(dp.rf._abc_6362_n9789) );
	NOR2X1 NOR2X1_1177 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9778), .B(dp.rf._abc_6362_n9789), .Y(dp.rf._abc_6362_n9790) );
	NOR2X1 NOR2X1_1178 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9790), .Y(dp.rf._abc_6362_n9791) );
	NAND2X1 NAND2X1_6607 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9768), .B(dp.rf._abc_6362_n9791), .Y(dp.rf._abc_6362_n9792) );
	NAND2X1 NAND2X1_6608 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n9792), .Y(dp.rf._abc_6362_n9793) );
	NOR2X1 NOR2X1_1179 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9746), .B(dp.rf._abc_6362_n9793), .Y(writedata_12__RAW) );
	NAND2X1 NAND2X1_6609 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<13>), .Y(dp.rf._abc_6362_n9795) );
	NAND2X1 NAND2X1_6610 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9795), .Y(dp.rf._abc_6362_n9796) );
	NOR2X1 NOR2X1_1180 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6670), .Y(dp.rf._abc_6362_n9797) );
	NOR2X1 NOR2X1_1181 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9796), .B(dp.rf._abc_6362_n9797), .Y(dp.rf._abc_6362_n9798) );
	NAND2X1 NAND2X1_6611 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<13>), .Y(dp.rf._abc_6362_n9799) );
	NAND2X1 NAND2X1_6612 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9799), .Y(dp.rf._abc_6362_n9800) );
	NOR2X1 NOR2X1_1182 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6675), .Y(dp.rf._abc_6362_n9801) );
	NOR2X1 NOR2X1_1183 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9800), .B(dp.rf._abc_6362_n9801), .Y(dp.rf._abc_6362_n9802) );
	NOR2X1 NOR2X1_1184 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9798), .B(dp.rf._abc_6362_n9802), .Y(dp.rf._abc_6362_n9803) );
	NAND2X1 NAND2X1_6613 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9803), .Y(dp.rf._abc_6362_n9804) );
	NAND2X1 NAND2X1_6614 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<13>), .Y(dp.rf._abc_6362_n9805) );
	NAND2X1 NAND2X1_6615 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9805), .Y(dp.rf._abc_6362_n9806) );
	NOR2X1 NOR2X1_1185 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6682), .Y(dp.rf._abc_6362_n9807) );
	NOR2X1 NOR2X1_1186 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9806), .B(dp.rf._abc_6362_n9807), .Y(dp.rf._abc_6362_n9808) );
	NAND2X1 NAND2X1_6616 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<13>), .Y(dp.rf._abc_6362_n9809) );
	NAND2X1 NAND2X1_6617 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9809), .Y(dp.rf._abc_6362_n9810) );
	NOR2X1 NOR2X1_1187 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6687), .Y(dp.rf._abc_6362_n9811) );
	NOR2X1 NOR2X1_1188 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9810), .B(dp.rf._abc_6362_n9811), .Y(dp.rf._abc_6362_n9812) );
	NOR2X1 NOR2X1_1189 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9808), .B(dp.rf._abc_6362_n9812), .Y(dp.rf._abc_6362_n9813) );
	NAND2X1 NAND2X1_6618 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9813), .Y(dp.rf._abc_6362_n9814) );
	NAND2X1 NAND2X1_6619 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9804), .B(dp.rf._abc_6362_n9814), .Y(dp.rf._abc_6362_n9815) );
	NAND2X1 NAND2X1_6620 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9815), .Y(dp.rf._abc_6362_n9816) );
	NAND2X1 NAND2X1_6621 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9816), .Y(dp.rf._abc_6362_n9817) );
	NAND2X1 NAND2X1_6622 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9818) );
	NOR2X1 NOR2X1_1190 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6696), .Y(dp.rf._abc_6362_n9819) );
	NOR2X1 NOR2X1_1191 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9819), .Y(dp.rf._abc_6362_n9820) );
	NAND2X1 NAND2X1_6623 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9818), .B(dp.rf._abc_6362_n9820), .Y(dp.rf._abc_6362_n9821) );
	NAND2X1 NAND2X1_6624 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9822) );
	NOR2X1 NOR2X1_1192 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6701), .Y(dp.rf._abc_6362_n9823) );
	NOR2X1 NOR2X1_1193 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9823), .Y(dp.rf._abc_6362_n9824) );
	NAND2X1 NAND2X1_6625 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9822), .B(dp.rf._abc_6362_n9824), .Y(dp.rf._abc_6362_n9825) );
	NAND2X1 NAND2X1_6626 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9821), .B(dp.rf._abc_6362_n9825), .Y(dp.rf._abc_6362_n9826) );
	NOR2X1 NOR2X1_1194 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9826), .Y(dp.rf._abc_6362_n9827) );
	NAND2X1 NAND2X1_6627 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9828) );
	NOR2X1 NOR2X1_1195 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6708), .Y(dp.rf._abc_6362_n9829) );
	NOR2X1 NOR2X1_1196 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9829), .Y(dp.rf._abc_6362_n9830) );
	NAND2X1 NAND2X1_6628 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9828), .B(dp.rf._abc_6362_n9830), .Y(dp.rf._abc_6362_n9831) );
	NAND2X1 NAND2X1_6629 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9832) );
	NOR2X1 NOR2X1_1197 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6713), .Y(dp.rf._abc_6362_n9833) );
	NOR2X1 NOR2X1_1198 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9833), .Y(dp.rf._abc_6362_n9834) );
	NAND2X1 NAND2X1_6630 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9832), .B(dp.rf._abc_6362_n9834), .Y(dp.rf._abc_6362_n9835) );
	NAND2X1 NAND2X1_6631 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9831), .B(dp.rf._abc_6362_n9835), .Y(dp.rf._abc_6362_n9836) );
	NOR2X1 NOR2X1_1199 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9836), .Y(dp.rf._abc_6362_n9837) );
	NOR2X1 NOR2X1_1200 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9827), .B(dp.rf._abc_6362_n9837), .Y(dp.rf._abc_6362_n9838) );
	NOR2X1 NOR2X1_1201 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9838), .Y(dp.rf._abc_6362_n9839) );
	NOR2X1 NOR2X1_1202 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9817), .B(dp.rf._abc_6362_n9839), .Y(dp.rf._abc_6362_n9840) );
	NAND2X1 NAND2X1_6632 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<13>), .Y(dp.rf._abc_6362_n9841) );
	NAND2X1 NAND2X1_6633 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9842) );
	NAND2X1 NAND2X1_6634 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9841), .B(dp.rf._abc_6362_n9842), .Y(dp.rf._abc_6362_n9843) );
	NAND2X1 NAND2X1_6635 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9843), .Y(dp.rf._abc_6362_n9844) );
	NAND2X1 NAND2X1_6636 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<13>), .Y(dp.rf._abc_6362_n9845) );
	NAND2X1 NAND2X1_6637 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9846) );
	NAND2X1 NAND2X1_6638 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9845), .B(dp.rf._abc_6362_n9846), .Y(dp.rf._abc_6362_n9847) );
	NAND2X1 NAND2X1_6639 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9847), .Y(dp.rf._abc_6362_n9848) );
	AND2X2 AND2X2_454 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9844), .B(dp.rf._abc_6362_n9848), .Y(dp.rf._abc_6362_n9849) );
	NAND2X1 NAND2X1_6640 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9849), .Y(dp.rf._abc_6362_n9850) );
	NAND2X1 NAND2X1_6641 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<13>), .Y(dp.rf._abc_6362_n9851) );
	NAND2X1 NAND2X1_6642 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9852) );
	NAND2X1 NAND2X1_6643 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9851), .B(dp.rf._abc_6362_n9852), .Y(dp.rf._abc_6362_n9853) );
	NAND2X1 NAND2X1_6644 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9853), .Y(dp.rf._abc_6362_n9854) );
	NAND2X1 NAND2X1_6645 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<13>), .Y(dp.rf._abc_6362_n9855) );
	NAND2X1 NAND2X1_6646 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9856) );
	NAND2X1 NAND2X1_6647 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9855), .B(dp.rf._abc_6362_n9856), .Y(dp.rf._abc_6362_n9857) );
	NAND2X1 NAND2X1_6648 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9857), .Y(dp.rf._abc_6362_n9858) );
	AND2X2 AND2X2_455 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9854), .B(dp.rf._abc_6362_n9858), .Y(dp.rf._abc_6362_n9859) );
	NAND2X1 NAND2X1_6649 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9859), .Y(dp.rf._abc_6362_n9860) );
	AND2X2 AND2X2_456 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9860), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n9861) );
	NAND2X1 NAND2X1_6650 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9850), .B(dp.rf._abc_6362_n9861), .Y(dp.rf._abc_6362_n9862) );
	NAND2X1 NAND2X1_6651 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9863) );
	NAND2X1 NAND2X1_6652 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<13>), .Y(dp.rf._abc_6362_n9864) );
	AND2X2 AND2X2_457 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9864), .B(instr[17]), .Y(dp.rf._abc_6362_n9865) );
	NAND2X1 NAND2X1_6653 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9863), .B(dp.rf._abc_6362_n9865), .Y(dp.rf._abc_6362_n9866) );
	NAND2X1 NAND2X1_6654 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9867) );
	NAND2X1 NAND2X1_6655 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<13>), .Y(dp.rf._abc_6362_n9868) );
	AND2X2 AND2X2_458 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9868), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9869) );
	NAND2X1 NAND2X1_6656 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9867), .B(dp.rf._abc_6362_n9869), .Y(dp.rf._abc_6362_n9870) );
	NAND2X1 NAND2X1_6657 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9866), .B(dp.rf._abc_6362_n9870), .Y(dp.rf._abc_6362_n9871) );
	AND2X2 AND2X2_459 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9871), .B(instr[18]), .Y(dp.rf._abc_6362_n9872) );
	NAND2X1 NAND2X1_6658 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9873) );
	NAND2X1 NAND2X1_6659 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<13>), .Y(dp.rf._abc_6362_n9874) );
	AND2X2 AND2X2_460 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9874), .B(instr[17]), .Y(dp.rf._abc_6362_n9875) );
	NAND2X1 NAND2X1_6660 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9873), .B(dp.rf._abc_6362_n9875), .Y(dp.rf._abc_6362_n9876) );
	NAND2X1 NAND2X1_6661 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<13>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9877) );
	NAND2X1 NAND2X1_6662 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<13>), .Y(dp.rf._abc_6362_n9878) );
	AND2X2 AND2X2_461 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9878), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9879) );
	NAND2X1 NAND2X1_6663 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9877), .B(dp.rf._abc_6362_n9879), .Y(dp.rf._abc_6362_n9880) );
	NAND2X1 NAND2X1_6664 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9876), .B(dp.rf._abc_6362_n9880), .Y(dp.rf._abc_6362_n9881) );
	NAND2X1 NAND2X1_6665 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9881), .Y(dp.rf._abc_6362_n9882) );
	NAND2X1 NAND2X1_6666 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9882), .Y(dp.rf._abc_6362_n9883) );
	NOR2X1 NOR2X1_1203 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9872), .B(dp.rf._abc_6362_n9883), .Y(dp.rf._abc_6362_n9884) );
	NOR2X1 NOR2X1_1204 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9884), .Y(dp.rf._abc_6362_n9885) );
	NAND2X1 NAND2X1_6667 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9862), .B(dp.rf._abc_6362_n9885), .Y(dp.rf._abc_6362_n9886) );
	NAND2X1 NAND2X1_6668 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n9886), .Y(dp.rf._abc_6362_n9887) );
	NOR2X1 NOR2X1_1205 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9840), .B(dp.rf._abc_6362_n9887), .Y(writedata_13__RAW) );
	NAND2X1 NAND2X1_6669 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<14>), .Y(dp.rf._abc_6362_n9889) );
	NAND2X1 NAND2X1_6670 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9889), .Y(dp.rf._abc_6362_n9890) );
	NOR2X1 NOR2X1_1206 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6772), .Y(dp.rf._abc_6362_n9891) );
	NOR2X1 NOR2X1_1207 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9890), .B(dp.rf._abc_6362_n9891), .Y(dp.rf._abc_6362_n9892) );
	NAND2X1 NAND2X1_6671 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<14>), .Y(dp.rf._abc_6362_n9893) );
	NAND2X1 NAND2X1_6672 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9893), .Y(dp.rf._abc_6362_n9894) );
	NOR2X1 NOR2X1_1208 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6777), .Y(dp.rf._abc_6362_n9895) );
	NOR2X1 NOR2X1_1209 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9894), .B(dp.rf._abc_6362_n9895), .Y(dp.rf._abc_6362_n9896) );
	NOR2X1 NOR2X1_1210 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9892), .B(dp.rf._abc_6362_n9896), .Y(dp.rf._abc_6362_n9897) );
	NAND2X1 NAND2X1_6673 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9897), .Y(dp.rf._abc_6362_n9898) );
	NAND2X1 NAND2X1_6674 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<14>), .Y(dp.rf._abc_6362_n9899) );
	NAND2X1 NAND2X1_6675 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9899), .Y(dp.rf._abc_6362_n9900) );
	NOR2X1 NOR2X1_1211 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6784), .Y(dp.rf._abc_6362_n9901) );
	NOR2X1 NOR2X1_1212 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9900), .B(dp.rf._abc_6362_n9901), .Y(dp.rf._abc_6362_n9902) );
	NAND2X1 NAND2X1_6676 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<14>), .Y(dp.rf._abc_6362_n9903) );
	NAND2X1 NAND2X1_6677 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9903), .Y(dp.rf._abc_6362_n9904) );
	NOR2X1 NOR2X1_1213 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n6789), .Y(dp.rf._abc_6362_n9905) );
	NOR2X1 NOR2X1_1214 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9904), .B(dp.rf._abc_6362_n9905), .Y(dp.rf._abc_6362_n9906) );
	NOR2X1 NOR2X1_1215 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9902), .B(dp.rf._abc_6362_n9906), .Y(dp.rf._abc_6362_n9907) );
	NAND2X1 NAND2X1_6678 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9907), .Y(dp.rf._abc_6362_n9908) );
	NAND2X1 NAND2X1_6679 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9898), .B(dp.rf._abc_6362_n9908), .Y(dp.rf._abc_6362_n9909) );
	NAND2X1 NAND2X1_6680 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9909), .Y(dp.rf._abc_6362_n9910) );
	NAND2X1 NAND2X1_6681 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9910), .Y(dp.rf._abc_6362_n9911) );
	NAND2X1 NAND2X1_6682 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9912) );
	NOR2X1 NOR2X1_1216 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6798), .Y(dp.rf._abc_6362_n9913) );
	NOR2X1 NOR2X1_1217 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9913), .Y(dp.rf._abc_6362_n9914) );
	NAND2X1 NAND2X1_6683 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9912), .B(dp.rf._abc_6362_n9914), .Y(dp.rf._abc_6362_n9915) );
	NAND2X1 NAND2X1_6684 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9916) );
	NOR2X1 NOR2X1_1218 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6803), .Y(dp.rf._abc_6362_n9917) );
	NOR2X1 NOR2X1_1219 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9917), .Y(dp.rf._abc_6362_n9918) );
	NAND2X1 NAND2X1_6685 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9916), .B(dp.rf._abc_6362_n9918), .Y(dp.rf._abc_6362_n9919) );
	NAND2X1 NAND2X1_6686 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9915), .B(dp.rf._abc_6362_n9919), .Y(dp.rf._abc_6362_n9920) );
	NOR2X1 NOR2X1_1220 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9920), .Y(dp.rf._abc_6362_n9921) );
	NAND2X1 NAND2X1_6687 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9922) );
	NOR2X1 NOR2X1_1221 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6810), .Y(dp.rf._abc_6362_n9923) );
	NOR2X1 NOR2X1_1222 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9923), .Y(dp.rf._abc_6362_n9924) );
	NAND2X1 NAND2X1_6688 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9922), .B(dp.rf._abc_6362_n9924), .Y(dp.rf._abc_6362_n9925) );
	NAND2X1 NAND2X1_6689 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9926) );
	NOR2X1 NOR2X1_1223 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n6815), .Y(dp.rf._abc_6362_n9927) );
	NOR2X1 NOR2X1_1224 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9927), .Y(dp.rf._abc_6362_n9928) );
	NAND2X1 NAND2X1_6690 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9926), .B(dp.rf._abc_6362_n9928), .Y(dp.rf._abc_6362_n9929) );
	NAND2X1 NAND2X1_6691 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9925), .B(dp.rf._abc_6362_n9929), .Y(dp.rf._abc_6362_n9930) );
	NOR2X1 NOR2X1_1225 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9930), .Y(dp.rf._abc_6362_n9931) );
	NOR2X1 NOR2X1_1226 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9921), .B(dp.rf._abc_6362_n9931), .Y(dp.rf._abc_6362_n9932) );
	NOR2X1 NOR2X1_1227 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n9932), .Y(dp.rf._abc_6362_n9933) );
	NOR2X1 NOR2X1_1228 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9911), .B(dp.rf._abc_6362_n9933), .Y(dp.rf._abc_6362_n9934) );
	NAND2X1 NAND2X1_6692 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<14>), .Y(dp.rf._abc_6362_n9935) );
	NAND2X1 NAND2X1_6693 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9936) );
	NAND2X1 NAND2X1_6694 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9935), .B(dp.rf._abc_6362_n9936), .Y(dp.rf._abc_6362_n9937) );
	NAND2X1 NAND2X1_6695 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9937), .Y(dp.rf._abc_6362_n9938) );
	NAND2X1 NAND2X1_6696 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<14>), .Y(dp.rf._abc_6362_n9939) );
	NAND2X1 NAND2X1_6697 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9940) );
	NAND2X1 NAND2X1_6698 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9939), .B(dp.rf._abc_6362_n9940), .Y(dp.rf._abc_6362_n9941) );
	NAND2X1 NAND2X1_6699 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9941), .Y(dp.rf._abc_6362_n9942) );
	AND2X2 AND2X2_462 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9938), .B(dp.rf._abc_6362_n9942), .Y(dp.rf._abc_6362_n9943) );
	NAND2X1 NAND2X1_6700 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9943), .Y(dp.rf._abc_6362_n9944) );
	NAND2X1 NAND2X1_6701 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<14>), .Y(dp.rf._abc_6362_n9945) );
	NAND2X1 NAND2X1_6702 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9946) );
	NAND2X1 NAND2X1_6703 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9945), .B(dp.rf._abc_6362_n9946), .Y(dp.rf._abc_6362_n9947) );
	NAND2X1 NAND2X1_6704 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9947), .Y(dp.rf._abc_6362_n9948) );
	NAND2X1 NAND2X1_6705 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<14>), .Y(dp.rf._abc_6362_n9949) );
	NAND2X1 NAND2X1_6706 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9950) );
	NAND2X1 NAND2X1_6707 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9949), .B(dp.rf._abc_6362_n9950), .Y(dp.rf._abc_6362_n9951) );
	NAND2X1 NAND2X1_6708 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9951), .Y(dp.rf._abc_6362_n9952) );
	AND2X2 AND2X2_463 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9948), .B(dp.rf._abc_6362_n9952), .Y(dp.rf._abc_6362_n9953) );
	NAND2X1 NAND2X1_6709 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9953), .Y(dp.rf._abc_6362_n9954) );
	AND2X2 AND2X2_464 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9954), .B(instr[19]), .Y(dp.rf._abc_6362_n9955) );
	NAND2X1 NAND2X1_6710 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9944), .B(dp.rf._abc_6362_n9955), .Y(dp.rf._abc_6362_n9956) );
	NAND2X1 NAND2X1_6711 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9957) );
	NAND2X1 NAND2X1_6712 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<14>), .Y(dp.rf._abc_6362_n9958) );
	AND2X2 AND2X2_465 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9958), .B(instr[17]), .Y(dp.rf._abc_6362_n9959) );
	NAND2X1 NAND2X1_6713 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9957), .B(dp.rf._abc_6362_n9959), .Y(dp.rf._abc_6362_n9960) );
	NAND2X1 NAND2X1_6714 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9961) );
	NAND2X1 NAND2X1_6715 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<14>), .Y(dp.rf._abc_6362_n9962) );
	AND2X2 AND2X2_466 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9962), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9963) );
	NAND2X1 NAND2X1_6716 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9961), .B(dp.rf._abc_6362_n9963), .Y(dp.rf._abc_6362_n9964) );
	NAND2X1 NAND2X1_6717 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9960), .B(dp.rf._abc_6362_n9964), .Y(dp.rf._abc_6362_n9965) );
	AND2X2 AND2X2_467 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9965), .B(instr[18]), .Y(dp.rf._abc_6362_n9966) );
	NAND2X1 NAND2X1_6718 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9967) );
	NAND2X1 NAND2X1_6719 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<14>), .Y(dp.rf._abc_6362_n9968) );
	AND2X2 AND2X2_468 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9968), .B(instr[17]), .Y(dp.rf._abc_6362_n9969) );
	NAND2X1 NAND2X1_6720 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9967), .B(dp.rf._abc_6362_n9969), .Y(dp.rf._abc_6362_n9970) );
	NAND2X1 NAND2X1_6721 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<14>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9971) );
	NAND2X1 NAND2X1_6722 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<14>), .Y(dp.rf._abc_6362_n9972) );
	AND2X2 AND2X2_469 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9972), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n9973) );
	NAND2X1 NAND2X1_6723 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9971), .B(dp.rf._abc_6362_n9973), .Y(dp.rf._abc_6362_n9974) );
	NAND2X1 NAND2X1_6724 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9970), .B(dp.rf._abc_6362_n9974), .Y(dp.rf._abc_6362_n9975) );
	NAND2X1 NAND2X1_6725 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n9975), .Y(dp.rf._abc_6362_n9976) );
	NAND2X1 NAND2X1_6726 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n9976), .Y(dp.rf._abc_6362_n9977) );
	NOR2X1 NOR2X1_1229 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9966), .B(dp.rf._abc_6362_n9977), .Y(dp.rf._abc_6362_n9978) );
	NOR2X1 NOR2X1_1230 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n9978), .Y(dp.rf._abc_6362_n9979) );
	NAND2X1 NAND2X1_6727 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9956), .B(dp.rf._abc_6362_n9979), .Y(dp.rf._abc_6362_n9980) );
	NAND2X1 NAND2X1_6728 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n9980), .Y(dp.rf._abc_6362_n9981) );
	NOR2X1 NOR2X1_1231 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9934), .B(dp.rf._abc_6362_n9981), .Y(writedata_14__RAW) );
	NAND2X1 NAND2X1_6729 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<15>), .Y(dp.rf._abc_6362_n9983) );
	NAND2X1 NAND2X1_6730 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9984) );
	NAND2X1 NAND2X1_6731 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9983), .B(dp.rf._abc_6362_n9984), .Y(dp.rf._abc_6362_n9985) );
	NAND2X1 NAND2X1_6732 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9985), .Y(dp.rf._abc_6362_n9986) );
	NAND2X1 NAND2X1_6733 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<15>), .Y(dp.rf._abc_6362_n9987) );
	NAND2X1 NAND2X1_6734 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9988) );
	NAND2X1 NAND2X1_6735 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9987), .B(dp.rf._abc_6362_n9988), .Y(dp.rf._abc_6362_n9989) );
	NAND2X1 NAND2X1_6736 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9989), .Y(dp.rf._abc_6362_n9990) );
	NAND2X1 NAND2X1_6737 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9986), .B(dp.rf._abc_6362_n9990), .Y(dp.rf._abc_6362_n9991) );
	NOR2X1 NOR2X1_1232 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n9991), .Y(dp.rf._abc_6362_n9992) );
	NAND2X1 NAND2X1_6738 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<15>), .Y(dp.rf._abc_6362_n9993) );
	NAND2X1 NAND2X1_6739 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9994) );
	NAND2X1 NAND2X1_6740 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9993), .B(dp.rf._abc_6362_n9994), .Y(dp.rf._abc_6362_n9995) );
	NAND2X1 NAND2X1_6741 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n9995), .Y(dp.rf._abc_6362_n9996) );
	NAND2X1 NAND2X1_6742 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<15>), .Y(dp.rf._abc_6362_n9997) );
	NAND2X1 NAND2X1_6743 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n9998) );
	NAND2X1 NAND2X1_6744 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9997), .B(dp.rf._abc_6362_n9998), .Y(dp.rf._abc_6362_n9999) );
	NAND2X1 NAND2X1_6745 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n9999), .Y(dp.rf._abc_6362_n10000) );
	AND2X2 AND2X2_470 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9996), .B(dp.rf._abc_6362_n10000), .Y(dp.rf._abc_6362_n10001) );
	NAND2X1 NAND2X1_6746 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10001), .Y(dp.rf._abc_6362_n10002) );
	NAND2X1 NAND2X1_6747 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10002), .Y(dp.rf._abc_6362_n10003) );
	NOR2X1 NOR2X1_1233 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n9992), .B(dp.rf._abc_6362_n10003), .Y(dp.rf._abc_6362_n10004) );
	NAND2X1 NAND2X1_6748 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<15>), .Y(dp.rf._abc_6362_n10005) );
	NAND2X1 NAND2X1_6749 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10006) );
	NAND2X1 NAND2X1_6750 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10005), .B(dp.rf._abc_6362_n10006), .Y(dp.rf._abc_6362_n10007) );
	NAND2X1 NAND2X1_6751 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10007), .Y(dp.rf._abc_6362_n10008) );
	NAND2X1 NAND2X1_6752 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<15>), .Y(dp.rf._abc_6362_n10009) );
	NAND2X1 NAND2X1_6753 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10010) );
	NAND2X1 NAND2X1_6754 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10009), .B(dp.rf._abc_6362_n10010), .Y(dp.rf._abc_6362_n10011) );
	NAND2X1 NAND2X1_6755 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10011), .Y(dp.rf._abc_6362_n10012) );
	AND2X2 AND2X2_471 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10008), .B(dp.rf._abc_6362_n10012), .Y(dp.rf._abc_6362_n10013) );
	NAND2X1 NAND2X1_6756 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10013), .Y(dp.rf._abc_6362_n10014) );
	NAND2X1 NAND2X1_6757 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<15>), .Y(dp.rf._abc_6362_n10015) );
	NAND2X1 NAND2X1_6758 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10015), .Y(dp.rf._abc_6362_n10016) );
	AND2X2 AND2X2_472 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf.rf_2_<15>), .Y(dp.rf._abc_6362_n10017) );
	NOR2X1 NOR2X1_1234 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10016), .B(dp.rf._abc_6362_n10017), .Y(dp.rf._abc_6362_n10018) );
	NAND2X1 NAND2X1_6759 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<15>), .Y(dp.rf._abc_6362_n10019) );
	NAND2X1 NAND2X1_6760 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10019), .Y(dp.rf._abc_6362_n10020) );
	INVX1 INVX1_257 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<15>), .Y(dp.rf._abc_6362_n10021) );
	NOR2X1 NOR2X1_1235 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n10021), .Y(dp.rf._abc_6362_n10022) );
	NOR2X1 NOR2X1_1236 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10020), .B(dp.rf._abc_6362_n10022), .Y(dp.rf._abc_6362_n10023) );
	OR2X2 OR2X2_103 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10018), .B(dp.rf._abc_6362_n10023), .Y(dp.rf._abc_6362_n10024) );
	NAND2X1 NAND2X1_6761 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10024), .Y(dp.rf._abc_6362_n10025) );
	AND2X2 AND2X2_473 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10025), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10026) );
	NAND2X1 NAND2X1_6762 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10014), .B(dp.rf._abc_6362_n10026), .Y(dp.rf._abc_6362_n10027) );
	NAND2X1 NAND2X1_6763 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10027), .Y(dp.rf._abc_6362_n10028) );
	NOR2X1 NOR2X1_1237 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10004), .B(dp.rf._abc_6362_n10028), .Y(dp.rf._abc_6362_n10029) );
	NAND2X1 NAND2X1_6764 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<15>), .Y(dp.rf._abc_6362_n10030) );
	NAND2X1 NAND2X1_6765 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10031) );
	NAND2X1 NAND2X1_6766 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10030), .B(dp.rf._abc_6362_n10031), .Y(dp.rf._abc_6362_n10032) );
	NAND2X1 NAND2X1_6767 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10032), .Y(dp.rf._abc_6362_n10033) );
	NAND2X1 NAND2X1_6768 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<15>), .Y(dp.rf._abc_6362_n10034) );
	NAND2X1 NAND2X1_6769 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10035) );
	NAND2X1 NAND2X1_6770 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10034), .B(dp.rf._abc_6362_n10035), .Y(dp.rf._abc_6362_n10036) );
	NAND2X1 NAND2X1_6771 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10036), .Y(dp.rf._abc_6362_n10037) );
	AND2X2 AND2X2_474 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10033), .B(dp.rf._abc_6362_n10037), .Y(dp.rf._abc_6362_n10038) );
	NAND2X1 NAND2X1_6772 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10038), .Y(dp.rf._abc_6362_n10039) );
	NAND2X1 NAND2X1_6773 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<15>), .Y(dp.rf._abc_6362_n10040) );
	NAND2X1 NAND2X1_6774 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10041) );
	NAND2X1 NAND2X1_6775 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10040), .B(dp.rf._abc_6362_n10041), .Y(dp.rf._abc_6362_n10042) );
	NAND2X1 NAND2X1_6776 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10042), .Y(dp.rf._abc_6362_n10043) );
	NAND2X1 NAND2X1_6777 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<15>), .Y(dp.rf._abc_6362_n10044) );
	NAND2X1 NAND2X1_6778 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10045) );
	NAND2X1 NAND2X1_6779 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10044), .B(dp.rf._abc_6362_n10045), .Y(dp.rf._abc_6362_n10046) );
	NAND2X1 NAND2X1_6780 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10046), .Y(dp.rf._abc_6362_n10047) );
	AND2X2 AND2X2_475 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10043), .B(dp.rf._abc_6362_n10047), .Y(dp.rf._abc_6362_n10048) );
	NAND2X1 NAND2X1_6781 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10048), .Y(dp.rf._abc_6362_n10049) );
	AND2X2 AND2X2_476 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10049), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10050) );
	NAND2X1 NAND2X1_6782 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10039), .B(dp.rf._abc_6362_n10050), .Y(dp.rf._abc_6362_n10051) );
	NAND2X1 NAND2X1_6783 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10052) );
	NAND2X1 NAND2X1_6784 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<15>), .Y(dp.rf._abc_6362_n10053) );
	AND2X2 AND2X2_477 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10053), .B(instr[17]), .Y(dp.rf._abc_6362_n10054) );
	NAND2X1 NAND2X1_6785 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10052), .B(dp.rf._abc_6362_n10054), .Y(dp.rf._abc_6362_n10055) );
	NAND2X1 NAND2X1_6786 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10056) );
	NAND2X1 NAND2X1_6787 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<15>), .Y(dp.rf._abc_6362_n10057) );
	AND2X2 AND2X2_478 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10057), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10058) );
	NAND2X1 NAND2X1_6788 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10056), .B(dp.rf._abc_6362_n10058), .Y(dp.rf._abc_6362_n10059) );
	NAND2X1 NAND2X1_6789 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10055), .B(dp.rf._abc_6362_n10059), .Y(dp.rf._abc_6362_n10060) );
	AND2X2 AND2X2_479 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10060), .B(instr[18]), .Y(dp.rf._abc_6362_n10061) );
	NAND2X1 NAND2X1_6790 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10062) );
	NAND2X1 NAND2X1_6791 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<15>), .Y(dp.rf._abc_6362_n10063) );
	AND2X2 AND2X2_480 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10063), .B(instr[17]), .Y(dp.rf._abc_6362_n10064) );
	NAND2X1 NAND2X1_6792 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10062), .B(dp.rf._abc_6362_n10064), .Y(dp.rf._abc_6362_n10065) );
	NAND2X1 NAND2X1_6793 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<15>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10066) );
	NAND2X1 NAND2X1_6794 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<15>), .Y(dp.rf._abc_6362_n10067) );
	AND2X2 AND2X2_481 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10067), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10068) );
	NAND2X1 NAND2X1_6795 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10066), .B(dp.rf._abc_6362_n10068), .Y(dp.rf._abc_6362_n10069) );
	NAND2X1 NAND2X1_6796 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10065), .B(dp.rf._abc_6362_n10069), .Y(dp.rf._abc_6362_n10070) );
	NAND2X1 NAND2X1_6797 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10070), .Y(dp.rf._abc_6362_n10071) );
	NAND2X1 NAND2X1_6798 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10071), .Y(dp.rf._abc_6362_n10072) );
	NOR2X1 NOR2X1_1238 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10061), .B(dp.rf._abc_6362_n10072), .Y(dp.rf._abc_6362_n10073) );
	NOR2X1 NOR2X1_1239 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10073), .Y(dp.rf._abc_6362_n10074) );
	NAND2X1 NAND2X1_6799 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10051), .B(dp.rf._abc_6362_n10074), .Y(dp.rf._abc_6362_n10075) );
	NAND2X1 NAND2X1_6800 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n10075), .Y(dp.rf._abc_6362_n10076) );
	NOR2X1 NOR2X1_1240 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10029), .B(dp.rf._abc_6362_n10076), .Y(writedata_15__RAW) );
	NAND2X1 NAND2X1_6801 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<16>), .Y(dp.rf._abc_6362_n10078) );
	NAND2X1 NAND2X1_6802 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10079) );
	NAND2X1 NAND2X1_6803 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10078), .B(dp.rf._abc_6362_n10079), .Y(dp.rf._abc_6362_n10080) );
	NAND2X1 NAND2X1_6804 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10080), .Y(dp.rf._abc_6362_n10081) );
	NAND2X1 NAND2X1_6805 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<16>), .Y(dp.rf._abc_6362_n10082) );
	NAND2X1 NAND2X1_6806 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10083) );
	NAND2X1 NAND2X1_6807 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10082), .B(dp.rf._abc_6362_n10083), .Y(dp.rf._abc_6362_n10084) );
	NAND2X1 NAND2X1_6808 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10084), .Y(dp.rf._abc_6362_n10085) );
	NAND2X1 NAND2X1_6809 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10081), .B(dp.rf._abc_6362_n10085), .Y(dp.rf._abc_6362_n10086) );
	NOR2X1 NOR2X1_1241 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10086), .Y(dp.rf._abc_6362_n10087) );
	NAND2X1 NAND2X1_6810 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<16>), .Y(dp.rf._abc_6362_n10088) );
	NAND2X1 NAND2X1_6811 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10089) );
	NAND2X1 NAND2X1_6812 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10088), .B(dp.rf._abc_6362_n10089), .Y(dp.rf._abc_6362_n10090) );
	NAND2X1 NAND2X1_6813 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10090), .Y(dp.rf._abc_6362_n10091) );
	NAND2X1 NAND2X1_6814 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<16>), .Y(dp.rf._abc_6362_n10092) );
	NAND2X1 NAND2X1_6815 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10093) );
	NAND2X1 NAND2X1_6816 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10092), .B(dp.rf._abc_6362_n10093), .Y(dp.rf._abc_6362_n10094) );
	NAND2X1 NAND2X1_6817 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10094), .Y(dp.rf._abc_6362_n10095) );
	AND2X2 AND2X2_482 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10091), .B(dp.rf._abc_6362_n10095), .Y(dp.rf._abc_6362_n10096) );
	NAND2X1 NAND2X1_6818 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10096), .Y(dp.rf._abc_6362_n10097) );
	NAND2X1 NAND2X1_6819 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n10097), .Y(dp.rf._abc_6362_n10098) );
	NOR2X1 NOR2X1_1242 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10087), .B(dp.rf._abc_6362_n10098), .Y(dp.rf._abc_6362_n10099) );
	NAND2X1 NAND2X1_6820 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<16>), .Y(dp.rf._abc_6362_n10100) );
	NAND2X1 NAND2X1_6821 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10101) );
	NAND2X1 NAND2X1_6822 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10100), .B(dp.rf._abc_6362_n10101), .Y(dp.rf._abc_6362_n10102) );
	NAND2X1 NAND2X1_6823 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10102), .Y(dp.rf._abc_6362_n10103) );
	NAND2X1 NAND2X1_6824 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<16>), .Y(dp.rf._abc_6362_n10104) );
	NAND2X1 NAND2X1_6825 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10105) );
	NAND2X1 NAND2X1_6826 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10104), .B(dp.rf._abc_6362_n10105), .Y(dp.rf._abc_6362_n10106) );
	NAND2X1 NAND2X1_6827 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10106), .Y(dp.rf._abc_6362_n10107) );
	NAND2X1 NAND2X1_6828 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10103), .B(dp.rf._abc_6362_n10107), .Y(dp.rf._abc_6362_n10108) );
	NAND2X1 NAND2X1_6829 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10108), .Y(dp.rf._abc_6362_n10109) );
	NAND2X1 NAND2X1_6830 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<16>), .Y(dp.rf._abc_6362_n10110) );
	NAND2X1 NAND2X1_6831 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10111) );
	NAND2X1 NAND2X1_6832 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10110), .B(dp.rf._abc_6362_n10111), .Y(dp.rf._abc_6362_n10112) );
	NAND2X1 NAND2X1_6833 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10112), .Y(dp.rf._abc_6362_n10113) );
	NAND2X1 NAND2X1_6834 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<16>), .Y(dp.rf._abc_6362_n10114) );
	NAND2X1 NAND2X1_6835 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10115) );
	NAND2X1 NAND2X1_6836 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10114), .B(dp.rf._abc_6362_n10115), .Y(dp.rf._abc_6362_n10116) );
	NAND2X1 NAND2X1_6837 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10116), .Y(dp.rf._abc_6362_n10117) );
	NAND2X1 NAND2X1_6838 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10113), .B(dp.rf._abc_6362_n10117), .Y(dp.rf._abc_6362_n10118) );
	NAND2X1 NAND2X1_6839 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10118), .Y(dp.rf._abc_6362_n10119) );
	NAND2X1 NAND2X1_6840 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10109), .B(dp.rf._abc_6362_n10119), .Y(dp.rf._abc_6362_n10120) );
	NAND2X1 NAND2X1_6841 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10120), .Y(dp.rf._abc_6362_n10121) );
	NAND2X1 NAND2X1_6842 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10121), .Y(dp.rf._abc_6362_n10122) );
	NOR2X1 NOR2X1_1243 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10099), .B(dp.rf._abc_6362_n10122), .Y(dp.rf._abc_6362_n10123) );
	NAND2X1 NAND2X1_6843 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<16>), .Y(dp.rf._abc_6362_n10124) );
	NAND2X1 NAND2X1_6844 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10124), .Y(dp.rf._abc_6362_n10125) );
	NOR2X1 NOR2X1_1244 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7016), .Y(dp.rf._abc_6362_n10126) );
	NOR2X1 NOR2X1_1245 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10125), .B(dp.rf._abc_6362_n10126), .Y(dp.rf._abc_6362_n10127) );
	NAND2X1 NAND2X1_6845 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<16>), .Y(dp.rf._abc_6362_n10128) );
	NAND2X1 NAND2X1_6846 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10128), .Y(dp.rf._abc_6362_n10129) );
	NOR2X1 NOR2X1_1246 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7021), .Y(dp.rf._abc_6362_n10130) );
	NOR2X1 NOR2X1_1247 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10129), .B(dp.rf._abc_6362_n10130), .Y(dp.rf._abc_6362_n10131) );
	OR2X2 OR2X2_104 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10127), .B(dp.rf._abc_6362_n10131), .Y(dp.rf._abc_6362_n10132) );
	NAND2X1 NAND2X1_6847 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10132), .Y(dp.rf._abc_6362_n10133) );
	NAND2X1 NAND2X1_6848 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<16>), .Y(dp.rf._abc_6362_n10134) );
	NAND2X1 NAND2X1_6849 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10134), .Y(dp.rf._abc_6362_n10135) );
	NOR2X1 NOR2X1_1248 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7028), .Y(dp.rf._abc_6362_n10136) );
	NOR2X1 NOR2X1_1249 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10135), .B(dp.rf._abc_6362_n10136), .Y(dp.rf._abc_6362_n10137) );
	NAND2X1 NAND2X1_6850 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<16>), .Y(dp.rf._abc_6362_n10138) );
	NAND2X1 NAND2X1_6851 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10138), .Y(dp.rf._abc_6362_n10139) );
	NOR2X1 NOR2X1_1250 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7033), .Y(dp.rf._abc_6362_n10140) );
	NOR2X1 NOR2X1_1251 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10139), .B(dp.rf._abc_6362_n10140), .Y(dp.rf._abc_6362_n10141) );
	OR2X2 OR2X2_105 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10137), .B(dp.rf._abc_6362_n10141), .Y(dp.rf._abc_6362_n10142) );
	NAND2X1 NAND2X1_6852 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10142), .Y(dp.rf._abc_6362_n10143) );
	AND2X2 AND2X2_483 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10143), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10144) );
	NAND2X1 NAND2X1_6853 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10133), .B(dp.rf._abc_6362_n10144), .Y(dp.rf._abc_6362_n10145) );
	NAND2X1 NAND2X1_6854 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10146) );
	NAND2X1 NAND2X1_6855 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<16>), .Y(dp.rf._abc_6362_n10147) );
	AND2X2 AND2X2_484 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10147), .B(instr[17]), .Y(dp.rf._abc_6362_n10148) );
	NAND2X1 NAND2X1_6856 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10146), .B(dp.rf._abc_6362_n10148), .Y(dp.rf._abc_6362_n10149) );
	NAND2X1 NAND2X1_6857 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10150) );
	NAND2X1 NAND2X1_6858 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<16>), .Y(dp.rf._abc_6362_n10151) );
	AND2X2 AND2X2_485 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10151), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10152) );
	NAND2X1 NAND2X1_6859 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10150), .B(dp.rf._abc_6362_n10152), .Y(dp.rf._abc_6362_n10153) );
	NAND2X1 NAND2X1_6860 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10149), .B(dp.rf._abc_6362_n10153), .Y(dp.rf._abc_6362_n10154) );
	AND2X2 AND2X2_486 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10154), .B(instr[18]), .Y(dp.rf._abc_6362_n10155) );
	NAND2X1 NAND2X1_6861 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10156) );
	NAND2X1 NAND2X1_6862 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<16>), .Y(dp.rf._abc_6362_n10157) );
	AND2X2 AND2X2_487 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10157), .B(instr[17]), .Y(dp.rf._abc_6362_n10158) );
	NAND2X1 NAND2X1_6863 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10156), .B(dp.rf._abc_6362_n10158), .Y(dp.rf._abc_6362_n10159) );
	NAND2X1 NAND2X1_6864 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<16>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10160) );
	NAND2X1 NAND2X1_6865 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<16>), .Y(dp.rf._abc_6362_n10161) );
	AND2X2 AND2X2_488 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10161), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10162) );
	NAND2X1 NAND2X1_6866 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10160), .B(dp.rf._abc_6362_n10162), .Y(dp.rf._abc_6362_n10163) );
	NAND2X1 NAND2X1_6867 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10159), .B(dp.rf._abc_6362_n10163), .Y(dp.rf._abc_6362_n10164) );
	NAND2X1 NAND2X1_6868 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10164), .Y(dp.rf._abc_6362_n10165) );
	NAND2X1 NAND2X1_6869 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10165), .Y(dp.rf._abc_6362_n10166) );
	NOR2X1 NOR2X1_1252 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10155), .B(dp.rf._abc_6362_n10166), .Y(dp.rf._abc_6362_n10167) );
	NOR2X1 NOR2X1_1253 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10167), .Y(dp.rf._abc_6362_n10168) );
	NAND2X1 NAND2X1_6870 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10145), .B(dp.rf._abc_6362_n10168), .Y(dp.rf._abc_6362_n10169) );
	NAND2X1 NAND2X1_6871 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n10169), .Y(dp.rf._abc_6362_n10170) );
	NOR2X1 NOR2X1_1254 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10123), .B(dp.rf._abc_6362_n10170), .Y(writedata_16__RAW) );
	NAND2X1 NAND2X1_6872 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<17>), .Y(dp.rf._abc_6362_n10172) );
	NAND2X1 NAND2X1_6873 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10172), .Y(dp.rf._abc_6362_n10173) );
	NOR2X1 NOR2X1_1255 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7090), .Y(dp.rf._abc_6362_n10174) );
	NOR2X1 NOR2X1_1256 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10173), .B(dp.rf._abc_6362_n10174), .Y(dp.rf._abc_6362_n10175) );
	NAND2X1 NAND2X1_6874 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<17>), .Y(dp.rf._abc_6362_n10176) );
	NAND2X1 NAND2X1_6875 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10176), .Y(dp.rf._abc_6362_n10177) );
	NOR2X1 NOR2X1_1257 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7095), .Y(dp.rf._abc_6362_n10178) );
	NOR2X1 NOR2X1_1258 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10177), .B(dp.rf._abc_6362_n10178), .Y(dp.rf._abc_6362_n10179) );
	NOR2X1 NOR2X1_1259 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10175), .B(dp.rf._abc_6362_n10179), .Y(dp.rf._abc_6362_n10180) );
	NAND2X1 NAND2X1_6876 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10180), .Y(dp.rf._abc_6362_n10181) );
	NAND2X1 NAND2X1_6877 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<17>), .Y(dp.rf._abc_6362_n10182) );
	NAND2X1 NAND2X1_6878 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10182), .Y(dp.rf._abc_6362_n10183) );
	NOR2X1 NOR2X1_1260 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7102), .Y(dp.rf._abc_6362_n10184) );
	NOR2X1 NOR2X1_1261 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10183), .B(dp.rf._abc_6362_n10184), .Y(dp.rf._abc_6362_n10185) );
	NAND2X1 NAND2X1_6879 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<17>), .Y(dp.rf._abc_6362_n10186) );
	NAND2X1 NAND2X1_6880 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10186), .Y(dp.rf._abc_6362_n10187) );
	NOR2X1 NOR2X1_1262 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7107), .Y(dp.rf._abc_6362_n10188) );
	NOR2X1 NOR2X1_1263 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10187), .B(dp.rf._abc_6362_n10188), .Y(dp.rf._abc_6362_n10189) );
	NOR2X1 NOR2X1_1264 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10185), .B(dp.rf._abc_6362_n10189), .Y(dp.rf._abc_6362_n10190) );
	NAND2X1 NAND2X1_6881 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10190), .Y(dp.rf._abc_6362_n10191) );
	NAND2X1 NAND2X1_6882 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10181), .B(dp.rf._abc_6362_n10191), .Y(dp.rf._abc_6362_n10192) );
	NAND2X1 NAND2X1_6883 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10192), .Y(dp.rf._abc_6362_n10193) );
	NAND2X1 NAND2X1_6884 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<17>), .Y(dp.rf._abc_6362_n10194) );
	NAND2X1 NAND2X1_6885 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<17>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10195) );
	NAND2X1 NAND2X1_6886 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10194), .B(dp.rf._abc_6362_n10195), .Y(dp.rf._abc_6362_n10196) );
	NAND2X1 NAND2X1_6887 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10196), .Y(dp.rf._abc_6362_n10197) );
	NAND2X1 NAND2X1_6888 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<17>), .Y(dp.rf._abc_6362_n10198) );
	NAND2X1 NAND2X1_6889 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<17>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10199) );
	NAND2X1 NAND2X1_6890 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10198), .B(dp.rf._abc_6362_n10199), .Y(dp.rf._abc_6362_n10200) );
	NAND2X1 NAND2X1_6891 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10200), .Y(dp.rf._abc_6362_n10201) );
	AND2X2 AND2X2_489 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10197), .B(dp.rf._abc_6362_n10201), .Y(dp.rf._abc_6362_n10202) );
	NAND2X1 NAND2X1_6892 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10202), .Y(dp.rf._abc_6362_n10203) );
	NAND2X1 NAND2X1_6893 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<17>), .Y(dp.rf._abc_6362_n10204) );
	NAND2X1 NAND2X1_6894 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10204), .Y(dp.rf._abc_6362_n10205) );
	AND2X2 AND2X2_490 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf.rf_2_<17>), .Y(dp.rf._abc_6362_n10206) );
	NOR2X1 NOR2X1_1265 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10205), .B(dp.rf._abc_6362_n10206), .Y(dp.rf._abc_6362_n10207) );
	NAND2X1 NAND2X1_6895 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<17>), .Y(dp.rf._abc_6362_n10208) );
	NAND2X1 NAND2X1_6896 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10208), .Y(dp.rf._abc_6362_n10209) );
	INVX1 INVX1_258 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<17>), .Y(dp.rf._abc_6362_n10210) );
	NOR2X1 NOR2X1_1266 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n10210), .Y(dp.rf._abc_6362_n10211) );
	NOR2X1 NOR2X1_1267 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10209), .B(dp.rf._abc_6362_n10211), .Y(dp.rf._abc_6362_n10212) );
	OR2X2 OR2X2_106 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10207), .B(dp.rf._abc_6362_n10212), .Y(dp.rf._abc_6362_n10213) );
	NAND2X1 NAND2X1_6897 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10213), .Y(dp.rf._abc_6362_n10214) );
	AND2X2 AND2X2_491 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10214), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10215) );
	NAND2X1 NAND2X1_6898 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10203), .B(dp.rf._abc_6362_n10215), .Y(dp.rf._abc_6362_n10216) );
	NAND2X1 NAND2X1_6899 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10193), .B(dp.rf._abc_6362_n10216), .Y(dp.rf._abc_6362_n10217) );
	NOR2X1 NOR2X1_1268 ( .gnd(gnd), .vdd(vdd), .A(instr[20]), .B(dp.rf._abc_6362_n10217), .Y(dp.rf._abc_6362_n10218) );
	NAND2X1 NAND2X1_6900 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<17>), .Y(dp.rf._abc_6362_n10219) );
	NAND2X1 NAND2X1_6901 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10219), .Y(dp.rf._abc_6362_n10220) );
	NOR2X1 NOR2X1_1269 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7118), .Y(dp.rf._abc_6362_n10221) );
	NOR2X1 NOR2X1_1270 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10220), .B(dp.rf._abc_6362_n10221), .Y(dp.rf._abc_6362_n10222) );
	NAND2X1 NAND2X1_6902 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<17>), .Y(dp.rf._abc_6362_n10223) );
	NAND2X1 NAND2X1_6903 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10223), .Y(dp.rf._abc_6362_n10224) );
	NOR2X1 NOR2X1_1271 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7123), .Y(dp.rf._abc_6362_n10225) );
	NOR2X1 NOR2X1_1272 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10224), .B(dp.rf._abc_6362_n10225), .Y(dp.rf._abc_6362_n10226) );
	OR2X2 OR2X2_107 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10222), .B(dp.rf._abc_6362_n10226), .Y(dp.rf._abc_6362_n10227) );
	NAND2X1 NAND2X1_6904 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10227), .Y(dp.rf._abc_6362_n10228) );
	NAND2X1 NAND2X1_6905 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<17>), .Y(dp.rf._abc_6362_n10229) );
	NAND2X1 NAND2X1_6906 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10229), .Y(dp.rf._abc_6362_n10230) );
	NOR2X1 NOR2X1_1273 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7130), .Y(dp.rf._abc_6362_n10231) );
	NOR2X1 NOR2X1_1274 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10230), .B(dp.rf._abc_6362_n10231), .Y(dp.rf._abc_6362_n10232) );
	NAND2X1 NAND2X1_6907 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<17>), .Y(dp.rf._abc_6362_n10233) );
	NAND2X1 NAND2X1_6908 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10233), .Y(dp.rf._abc_6362_n10234) );
	NOR2X1 NOR2X1_1275 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7135), .Y(dp.rf._abc_6362_n10235) );
	NOR2X1 NOR2X1_1276 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10234), .B(dp.rf._abc_6362_n10235), .Y(dp.rf._abc_6362_n10236) );
	OR2X2 OR2X2_108 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10232), .B(dp.rf._abc_6362_n10236), .Y(dp.rf._abc_6362_n10237) );
	NAND2X1 NAND2X1_6909 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10237), .Y(dp.rf._abc_6362_n10238) );
	AND2X2 AND2X2_492 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10238), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10239) );
	NAND2X1 NAND2X1_6910 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10228), .B(dp.rf._abc_6362_n10239), .Y(dp.rf._abc_6362_n10240) );
	NAND2X1 NAND2X1_6911 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<17>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10241) );
	NAND2X1 NAND2X1_6912 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<17>), .Y(dp.rf._abc_6362_n10242) );
	AND2X2 AND2X2_493 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10242), .B(instr[17]), .Y(dp.rf._abc_6362_n10243) );
	NAND2X1 NAND2X1_6913 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10241), .B(dp.rf._abc_6362_n10243), .Y(dp.rf._abc_6362_n10244) );
	NAND2X1 NAND2X1_6914 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<17>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10245) );
	NAND2X1 NAND2X1_6915 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<17>), .Y(dp.rf._abc_6362_n10246) );
	AND2X2 AND2X2_494 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10246), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10247) );
	NAND2X1 NAND2X1_6916 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10245), .B(dp.rf._abc_6362_n10247), .Y(dp.rf._abc_6362_n10248) );
	NAND2X1 NAND2X1_6917 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10244), .B(dp.rf._abc_6362_n10248), .Y(dp.rf._abc_6362_n10249) );
	AND2X2 AND2X2_495 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10249), .B(instr[18]), .Y(dp.rf._abc_6362_n10250) );
	NAND2X1 NAND2X1_6918 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<17>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10251) );
	NAND2X1 NAND2X1_6919 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<17>), .Y(dp.rf._abc_6362_n10252) );
	AND2X2 AND2X2_496 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10252), .B(instr[17]), .Y(dp.rf._abc_6362_n10253) );
	NAND2X1 NAND2X1_6920 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10251), .B(dp.rf._abc_6362_n10253), .Y(dp.rf._abc_6362_n10254) );
	NAND2X1 NAND2X1_6921 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<17>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10255) );
	NAND2X1 NAND2X1_6922 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<17>), .Y(dp.rf._abc_6362_n10256) );
	AND2X2 AND2X2_497 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10256), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10257) );
	NAND2X1 NAND2X1_6923 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10255), .B(dp.rf._abc_6362_n10257), .Y(dp.rf._abc_6362_n10258) );
	NAND2X1 NAND2X1_6924 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10254), .B(dp.rf._abc_6362_n10258), .Y(dp.rf._abc_6362_n10259) );
	NAND2X1 NAND2X1_6925 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10259), .Y(dp.rf._abc_6362_n10260) );
	NAND2X1 NAND2X1_6926 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10260), .Y(dp.rf._abc_6362_n10261) );
	NOR2X1 NOR2X1_1277 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10250), .B(dp.rf._abc_6362_n10261), .Y(dp.rf._abc_6362_n10262) );
	NOR2X1 NOR2X1_1278 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10262), .Y(dp.rf._abc_6362_n10263) );
	NAND2X1 NAND2X1_6927 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10240), .B(dp.rf._abc_6362_n10263), .Y(dp.rf._abc_6362_n10264) );
	NAND2X1 NAND2X1_6928 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n10264), .Y(dp.rf._abc_6362_n10265) );
	NOR2X1 NOR2X1_1279 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10218), .B(dp.rf._abc_6362_n10265), .Y(writedata_17__RAW) );
	NAND2X1 NAND2X1_6929 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<18>), .Y(dp.rf._abc_6362_n10267) );
	NAND2X1 NAND2X1_6930 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<18>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10268) );
	NAND2X1 NAND2X1_6931 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10267), .B(dp.rf._abc_6362_n10268), .Y(dp.rf._abc_6362_n10269) );
	NAND2X1 NAND2X1_6932 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10269), .Y(dp.rf._abc_6362_n10270) );
	NAND2X1 NAND2X1_6933 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<18>), .Y(dp.rf._abc_6362_n10271) );
	NAND2X1 NAND2X1_6934 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<18>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10272) );
	NAND2X1 NAND2X1_6935 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10271), .B(dp.rf._abc_6362_n10272), .Y(dp.rf._abc_6362_n10273) );
	NAND2X1 NAND2X1_6936 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10273), .Y(dp.rf._abc_6362_n10274) );
	NAND2X1 NAND2X1_6937 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10270), .B(dp.rf._abc_6362_n10274), .Y(dp.rf._abc_6362_n10275) );
	NOR2X1 NOR2X1_1280 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10275), .Y(dp.rf._abc_6362_n10276) );
	NAND2X1 NAND2X1_6938 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<18>), .Y(dp.rf._abc_6362_n10277) );
	NAND2X1 NAND2X1_6939 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<18>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10278) );
	NAND2X1 NAND2X1_6940 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10277), .B(dp.rf._abc_6362_n10278), .Y(dp.rf._abc_6362_n10279) );
	NAND2X1 NAND2X1_6941 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10279), .Y(dp.rf._abc_6362_n10280) );
	NAND2X1 NAND2X1_6942 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<18>), .Y(dp.rf._abc_6362_n10281) );
	NAND2X1 NAND2X1_6943 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<18>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10282) );
	NAND2X1 NAND2X1_6944 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10281), .B(dp.rf._abc_6362_n10282), .Y(dp.rf._abc_6362_n10283) );
	NAND2X1 NAND2X1_6945 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10283), .Y(dp.rf._abc_6362_n10284) );
	AND2X2 AND2X2_498 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10280), .B(dp.rf._abc_6362_n10284), .Y(dp.rf._abc_6362_n10285) );
	NAND2X1 NAND2X1_6946 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10285), .Y(dp.rf._abc_6362_n10286) );
	NAND2X1 NAND2X1_6947 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n10286), .Y(dp.rf._abc_6362_n10287) );
	NOR2X1 NOR2X1_1281 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10276), .B(dp.rf._abc_6362_n10287), .Y(dp.rf._abc_6362_n10288) );
	NAND2X1 NAND2X1_6948 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<18>), .Y(dp.rf._abc_6362_n10289) );
	NAND2X1 NAND2X1_6949 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10289), .Y(dp.rf._abc_6362_n10290) );
	NOR2X1 NOR2X1_1282 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7170), .Y(dp.rf._abc_6362_n10291) );
	NOR2X1 NOR2X1_1283 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10290), .B(dp.rf._abc_6362_n10291), .Y(dp.rf._abc_6362_n10292) );
	NAND2X1 NAND2X1_6950 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<18>), .Y(dp.rf._abc_6362_n10293) );
	NAND2X1 NAND2X1_6951 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10293), .Y(dp.rf._abc_6362_n10294) );
	NOR2X1 NOR2X1_1284 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7175), .Y(dp.rf._abc_6362_n10295) );
	NOR2X1 NOR2X1_1285 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10294), .B(dp.rf._abc_6362_n10295), .Y(dp.rf._abc_6362_n10296) );
	NOR2X1 NOR2X1_1286 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10292), .B(dp.rf._abc_6362_n10296), .Y(dp.rf._abc_6362_n10297) );
	NAND2X1 NAND2X1_6952 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10297), .Y(dp.rf._abc_6362_n10298) );
	NAND2X1 NAND2X1_6953 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<18>), .Y(dp.rf._abc_6362_n10299) );
	NAND2X1 NAND2X1_6954 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10299), .Y(dp.rf._abc_6362_n10300) );
	NOR2X1 NOR2X1_1287 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7182), .Y(dp.rf._abc_6362_n10301) );
	NOR2X1 NOR2X1_1288 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10300), .B(dp.rf._abc_6362_n10301), .Y(dp.rf._abc_6362_n10302) );
	NAND2X1 NAND2X1_6955 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<18>), .Y(dp.rf._abc_6362_n10303) );
	NAND2X1 NAND2X1_6956 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10303), .Y(dp.rf._abc_6362_n10304) );
	NOR2X1 NOR2X1_1289 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7187), .Y(dp.rf._abc_6362_n10305) );
	NOR2X1 NOR2X1_1290 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10304), .B(dp.rf._abc_6362_n10305), .Y(dp.rf._abc_6362_n10306) );
	NOR2X1 NOR2X1_1291 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10302), .B(dp.rf._abc_6362_n10306), .Y(dp.rf._abc_6362_n10307) );
	NAND2X1 NAND2X1_6957 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10307), .Y(dp.rf._abc_6362_n10308) );
	NAND2X1 NAND2X1_6958 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10298), .B(dp.rf._abc_6362_n10308), .Y(dp.rf._abc_6362_n10309) );
	NAND2X1 NAND2X1_6959 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10309), .Y(dp.rf._abc_6362_n10310) );
	NAND2X1 NAND2X1_6960 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10310), .Y(dp.rf._abc_6362_n10311) );
	NOR2X1 NOR2X1_1292 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10288), .B(dp.rf._abc_6362_n10311), .Y(dp.rf._abc_6362_n10312) );
	NAND2X1 NAND2X1_6961 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<18>), .Y(dp.rf._abc_6362_n10313) );
	NAND2X1 NAND2X1_6962 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10313), .Y(dp.rf._abc_6362_n10314) );
	NOR2X1 NOR2X1_1293 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7221), .Y(dp.rf._abc_6362_n10315) );
	NOR2X1 NOR2X1_1294 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10314), .B(dp.rf._abc_6362_n10315), .Y(dp.rf._abc_6362_n10316) );
	NAND2X1 NAND2X1_6963 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<18>), .Y(dp.rf._abc_6362_n10317) );
	NAND2X1 NAND2X1_6964 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10317), .Y(dp.rf._abc_6362_n10318) );
	NOR2X1 NOR2X1_1295 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7226), .Y(dp.rf._abc_6362_n10319) );
	NOR2X1 NOR2X1_1296 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10318), .B(dp.rf._abc_6362_n10319), .Y(dp.rf._abc_6362_n10320) );
	OR2X2 OR2X2_109 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10316), .B(dp.rf._abc_6362_n10320), .Y(dp.rf._abc_6362_n10321) );
	NAND2X1 NAND2X1_6965 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10321), .Y(dp.rf._abc_6362_n10322) );
	NAND2X1 NAND2X1_6966 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<18>), .Y(dp.rf._abc_6362_n10323) );
	NAND2X1 NAND2X1_6967 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10323), .Y(dp.rf._abc_6362_n10324) );
	NOR2X1 NOR2X1_1297 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7233), .Y(dp.rf._abc_6362_n10325) );
	NOR2X1 NOR2X1_1298 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10324), .B(dp.rf._abc_6362_n10325), .Y(dp.rf._abc_6362_n10326) );
	NAND2X1 NAND2X1_6968 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<18>), .Y(dp.rf._abc_6362_n10327) );
	NAND2X1 NAND2X1_6969 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10327), .Y(dp.rf._abc_6362_n10328) );
	NOR2X1 NOR2X1_1299 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7238), .Y(dp.rf._abc_6362_n10329) );
	NOR2X1 NOR2X1_1300 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10328), .B(dp.rf._abc_6362_n10329), .Y(dp.rf._abc_6362_n10330) );
	OR2X2 OR2X2_110 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10326), .B(dp.rf._abc_6362_n10330), .Y(dp.rf._abc_6362_n10331) );
	NAND2X1 NAND2X1_6970 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10331), .Y(dp.rf._abc_6362_n10332) );
	AND2X2 AND2X2_499 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10332), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10333) );
	NAND2X1 NAND2X1_6971 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10322), .B(dp.rf._abc_6362_n10333), .Y(dp.rf._abc_6362_n10334) );
	NAND2X1 NAND2X1_6972 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<18>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10335) );
	NAND2X1 NAND2X1_6973 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<18>), .Y(dp.rf._abc_6362_n10336) );
	AND2X2 AND2X2_500 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10336), .B(instr[17]), .Y(dp.rf._abc_6362_n10337) );
	NAND2X1 NAND2X1_6974 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10335), .B(dp.rf._abc_6362_n10337), .Y(dp.rf._abc_6362_n10338) );
	NAND2X1 NAND2X1_6975 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<18>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10339) );
	NAND2X1 NAND2X1_6976 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<18>), .Y(dp.rf._abc_6362_n10340) );
	AND2X2 AND2X2_501 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10340), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10341) );
	NAND2X1 NAND2X1_6977 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10339), .B(dp.rf._abc_6362_n10341), .Y(dp.rf._abc_6362_n10342) );
	NAND2X1 NAND2X1_6978 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10338), .B(dp.rf._abc_6362_n10342), .Y(dp.rf._abc_6362_n10343) );
	AND2X2 AND2X2_502 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10343), .B(instr[18]), .Y(dp.rf._abc_6362_n10344) );
	NAND2X1 NAND2X1_6979 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<18>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10345) );
	NAND2X1 NAND2X1_6980 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<18>), .Y(dp.rf._abc_6362_n10346) );
	AND2X2 AND2X2_503 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10346), .B(instr[17]), .Y(dp.rf._abc_6362_n10347) );
	NAND2X1 NAND2X1_6981 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10345), .B(dp.rf._abc_6362_n10347), .Y(dp.rf._abc_6362_n10348) );
	NAND2X1 NAND2X1_6982 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<18>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10349) );
	NAND2X1 NAND2X1_6983 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<18>), .Y(dp.rf._abc_6362_n10350) );
	AND2X2 AND2X2_504 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10350), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10351) );
	NAND2X1 NAND2X1_6984 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10349), .B(dp.rf._abc_6362_n10351), .Y(dp.rf._abc_6362_n10352) );
	NAND2X1 NAND2X1_6985 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10348), .B(dp.rf._abc_6362_n10352), .Y(dp.rf._abc_6362_n10353) );
	NAND2X1 NAND2X1_6986 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10353), .Y(dp.rf._abc_6362_n10354) );
	NAND2X1 NAND2X1_6987 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10354), .Y(dp.rf._abc_6362_n10355) );
	NOR2X1 NOR2X1_1301 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10344), .B(dp.rf._abc_6362_n10355), .Y(dp.rf._abc_6362_n10356) );
	NOR2X1 NOR2X1_1302 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10356), .Y(dp.rf._abc_6362_n10357) );
	NAND2X1 NAND2X1_6988 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10334), .B(dp.rf._abc_6362_n10357), .Y(dp.rf._abc_6362_n10358) );
	NAND2X1 NAND2X1_6989 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n10358), .Y(dp.rf._abc_6362_n10359) );
	NOR2X1 NOR2X1_1303 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10312), .B(dp.rf._abc_6362_n10359), .Y(writedata_18__RAW) );
	NAND2X1 NAND2X1_6990 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<19>), .Y(dp.rf._abc_6362_n10361) );
	NAND2X1 NAND2X1_6991 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10362) );
	NAND2X1 NAND2X1_6992 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10361), .B(dp.rf._abc_6362_n10362), .Y(dp.rf._abc_6362_n10363) );
	NAND2X1 NAND2X1_6993 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10363), .Y(dp.rf._abc_6362_n10364) );
	NAND2X1 NAND2X1_6994 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<19>), .Y(dp.rf._abc_6362_n10365) );
	NAND2X1 NAND2X1_6995 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10366) );
	NAND2X1 NAND2X1_6996 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10365), .B(dp.rf._abc_6362_n10366), .Y(dp.rf._abc_6362_n10367) );
	NAND2X1 NAND2X1_6997 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10367), .Y(dp.rf._abc_6362_n10368) );
	NAND2X1 NAND2X1_6998 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10364), .B(dp.rf._abc_6362_n10368), .Y(dp.rf._abc_6362_n10369) );
	NOR2X1 NOR2X1_1304 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10369), .Y(dp.rf._abc_6362_n10370) );
	NAND2X1 NAND2X1_6999 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<19>), .Y(dp.rf._abc_6362_n10371) );
	NAND2X1 NAND2X1_7000 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10372) );
	NAND2X1 NAND2X1_7001 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10371), .B(dp.rf._abc_6362_n10372), .Y(dp.rf._abc_6362_n10373) );
	NAND2X1 NAND2X1_7002 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10373), .Y(dp.rf._abc_6362_n10374) );
	NAND2X1 NAND2X1_7003 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<19>), .Y(dp.rf._abc_6362_n10375) );
	NAND2X1 NAND2X1_7004 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10376) );
	NAND2X1 NAND2X1_7005 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10375), .B(dp.rf._abc_6362_n10376), .Y(dp.rf._abc_6362_n10377) );
	NAND2X1 NAND2X1_7006 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10377), .Y(dp.rf._abc_6362_n10378) );
	AND2X2 AND2X2_505 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10374), .B(dp.rf._abc_6362_n10378), .Y(dp.rf._abc_6362_n10379) );
	NAND2X1 NAND2X1_7007 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10379), .Y(dp.rf._abc_6362_n10380) );
	NAND2X1 NAND2X1_7008 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10380), .Y(dp.rf._abc_6362_n10381) );
	NOR2X1 NOR2X1_1305 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10370), .B(dp.rf._abc_6362_n10381), .Y(dp.rf._abc_6362_n10382) );
	NAND2X1 NAND2X1_7009 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<19>), .Y(dp.rf._abc_6362_n10383) );
	NAND2X1 NAND2X1_7010 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10384) );
	NAND2X1 NAND2X1_7011 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10383), .B(dp.rf._abc_6362_n10384), .Y(dp.rf._abc_6362_n10385) );
	NAND2X1 NAND2X1_7012 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10385), .Y(dp.rf._abc_6362_n10386) );
	NAND2X1 NAND2X1_7013 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<19>), .Y(dp.rf._abc_6362_n10387) );
	NAND2X1 NAND2X1_7014 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10388) );
	NAND2X1 NAND2X1_7015 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10387), .B(dp.rf._abc_6362_n10388), .Y(dp.rf._abc_6362_n10389) );
	NAND2X1 NAND2X1_7016 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10389), .Y(dp.rf._abc_6362_n10390) );
	AND2X2 AND2X2_506 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10386), .B(dp.rf._abc_6362_n10390), .Y(dp.rf._abc_6362_n10391) );
	NAND2X1 NAND2X1_7017 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10391), .Y(dp.rf._abc_6362_n10392) );
	NAND2X1 NAND2X1_7018 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<19>), .Y(dp.rf._abc_6362_n10393) );
	NAND2X1 NAND2X1_7019 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10393), .Y(dp.rf._abc_6362_n10394) );
	AND2X2 AND2X2_507 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf.rf_2_<19>), .Y(dp.rf._abc_6362_n10395) );
	NOR2X1 NOR2X1_1306 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10394), .B(dp.rf._abc_6362_n10395), .Y(dp.rf._abc_6362_n10396) );
	NAND2X1 NAND2X1_7020 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<19>), .Y(dp.rf._abc_6362_n10397) );
	NAND2X1 NAND2X1_7021 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10397), .Y(dp.rf._abc_6362_n10398) );
	INVX1 INVX1_259 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<19>), .Y(dp.rf._abc_6362_n10399) );
	NOR2X1 NOR2X1_1307 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n10399), .Y(dp.rf._abc_6362_n10400) );
	NOR2X1 NOR2X1_1308 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10398), .B(dp.rf._abc_6362_n10400), .Y(dp.rf._abc_6362_n10401) );
	OR2X2 OR2X2_111 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10396), .B(dp.rf._abc_6362_n10401), .Y(dp.rf._abc_6362_n10402) );
	NAND2X1 NAND2X1_7022 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10402), .Y(dp.rf._abc_6362_n10403) );
	AND2X2 AND2X2_508 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10403), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10404) );
	NAND2X1 NAND2X1_7023 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10392), .B(dp.rf._abc_6362_n10404), .Y(dp.rf._abc_6362_n10405) );
	NAND2X1 NAND2X1_7024 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10405), .Y(dp.rf._abc_6362_n10406) );
	NOR2X1 NOR2X1_1309 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10382), .B(dp.rf._abc_6362_n10406), .Y(dp.rf._abc_6362_n10407) );
	NAND2X1 NAND2X1_7025 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<19>), .Y(dp.rf._abc_6362_n10408) );
	NAND2X1 NAND2X1_7026 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10409) );
	NAND2X1 NAND2X1_7027 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10408), .B(dp.rf._abc_6362_n10409), .Y(dp.rf._abc_6362_n10410) );
	NAND2X1 NAND2X1_7028 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10410), .Y(dp.rf._abc_6362_n10411) );
	NAND2X1 NAND2X1_7029 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<19>), .Y(dp.rf._abc_6362_n10412) );
	NAND2X1 NAND2X1_7030 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10413) );
	NAND2X1 NAND2X1_7031 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10412), .B(dp.rf._abc_6362_n10413), .Y(dp.rf._abc_6362_n10414) );
	NAND2X1 NAND2X1_7032 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10414), .Y(dp.rf._abc_6362_n10415) );
	AND2X2 AND2X2_509 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10411), .B(dp.rf._abc_6362_n10415), .Y(dp.rf._abc_6362_n10416) );
	NAND2X1 NAND2X1_7033 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10416), .Y(dp.rf._abc_6362_n10417) );
	NAND2X1 NAND2X1_7034 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<19>), .Y(dp.rf._abc_6362_n10418) );
	NAND2X1 NAND2X1_7035 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10419) );
	NAND2X1 NAND2X1_7036 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10418), .B(dp.rf._abc_6362_n10419), .Y(dp.rf._abc_6362_n10420) );
	NAND2X1 NAND2X1_7037 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10420), .Y(dp.rf._abc_6362_n10421) );
	NAND2X1 NAND2X1_7038 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<19>), .Y(dp.rf._abc_6362_n10422) );
	NAND2X1 NAND2X1_7039 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10423) );
	NAND2X1 NAND2X1_7040 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10422), .B(dp.rf._abc_6362_n10423), .Y(dp.rf._abc_6362_n10424) );
	NAND2X1 NAND2X1_7041 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10424), .Y(dp.rf._abc_6362_n10425) );
	AND2X2 AND2X2_510 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10421), .B(dp.rf._abc_6362_n10425), .Y(dp.rf._abc_6362_n10426) );
	NAND2X1 NAND2X1_7042 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10426), .Y(dp.rf._abc_6362_n10427) );
	AND2X2 AND2X2_511 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10427), .B(instr[19]), .Y(dp.rf._abc_6362_n10428) );
	NAND2X1 NAND2X1_7043 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10417), .B(dp.rf._abc_6362_n10428), .Y(dp.rf._abc_6362_n10429) );
	NAND2X1 NAND2X1_7044 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10430) );
	NAND2X1 NAND2X1_7045 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<19>), .Y(dp.rf._abc_6362_n10431) );
	AND2X2 AND2X2_512 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10431), .B(instr[17]), .Y(dp.rf._abc_6362_n10432) );
	NAND2X1 NAND2X1_7046 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10430), .B(dp.rf._abc_6362_n10432), .Y(dp.rf._abc_6362_n10433) );
	NAND2X1 NAND2X1_7047 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10434) );
	NAND2X1 NAND2X1_7048 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<19>), .Y(dp.rf._abc_6362_n10435) );
	AND2X2 AND2X2_513 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10435), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10436) );
	NAND2X1 NAND2X1_7049 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10434), .B(dp.rf._abc_6362_n10436), .Y(dp.rf._abc_6362_n10437) );
	NAND2X1 NAND2X1_7050 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10433), .B(dp.rf._abc_6362_n10437), .Y(dp.rf._abc_6362_n10438) );
	AND2X2 AND2X2_514 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10438), .B(instr[18]), .Y(dp.rf._abc_6362_n10439) );
	NAND2X1 NAND2X1_7051 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10440) );
	NAND2X1 NAND2X1_7052 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<19>), .Y(dp.rf._abc_6362_n10441) );
	AND2X2 AND2X2_515 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10441), .B(instr[17]), .Y(dp.rf._abc_6362_n10442) );
	NAND2X1 NAND2X1_7053 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10440), .B(dp.rf._abc_6362_n10442), .Y(dp.rf._abc_6362_n10443) );
	NAND2X1 NAND2X1_7054 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<19>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10444) );
	NAND2X1 NAND2X1_7055 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<19>), .Y(dp.rf._abc_6362_n10445) );
	AND2X2 AND2X2_516 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10445), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10446) );
	NAND2X1 NAND2X1_7056 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10444), .B(dp.rf._abc_6362_n10446), .Y(dp.rf._abc_6362_n10447) );
	NAND2X1 NAND2X1_7057 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10443), .B(dp.rf._abc_6362_n10447), .Y(dp.rf._abc_6362_n10448) );
	NAND2X1 NAND2X1_7058 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10448), .Y(dp.rf._abc_6362_n10449) );
	NAND2X1 NAND2X1_7059 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n10449), .Y(dp.rf._abc_6362_n10450) );
	NOR2X1 NOR2X1_1310 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10439), .B(dp.rf._abc_6362_n10450), .Y(dp.rf._abc_6362_n10451) );
	NOR2X1 NOR2X1_1311 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10451), .Y(dp.rf._abc_6362_n10452) );
	NAND2X1 NAND2X1_7060 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10429), .B(dp.rf._abc_6362_n10452), .Y(dp.rf._abc_6362_n10453) );
	NAND2X1 NAND2X1_7061 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n10453), .Y(dp.rf._abc_6362_n10454) );
	NOR2X1 NOR2X1_1312 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10407), .B(dp.rf._abc_6362_n10454), .Y(writedata_19__RAW) );
	NAND2X1 NAND2X1_7062 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<20>), .Y(dp.rf._abc_6362_n10456) );
	NAND2X1 NAND2X1_7063 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10457) );
	NAND2X1 NAND2X1_7064 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10456), .B(dp.rf._abc_6362_n10457), .Y(dp.rf._abc_6362_n10458) );
	NAND2X1 NAND2X1_7065 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10458), .Y(dp.rf._abc_6362_n10459) );
	NAND2X1 NAND2X1_7066 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<20>), .Y(dp.rf._abc_6362_n10460) );
	NAND2X1 NAND2X1_7067 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10461) );
	NAND2X1 NAND2X1_7068 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10460), .B(dp.rf._abc_6362_n10461), .Y(dp.rf._abc_6362_n10462) );
	NAND2X1 NAND2X1_7069 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10462), .Y(dp.rf._abc_6362_n10463) );
	NAND2X1 NAND2X1_7070 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10459), .B(dp.rf._abc_6362_n10463), .Y(dp.rf._abc_6362_n10464) );
	NOR2X1 NOR2X1_1313 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10464), .Y(dp.rf._abc_6362_n10465) );
	NAND2X1 NAND2X1_7071 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<20>), .Y(dp.rf._abc_6362_n10466) );
	NAND2X1 NAND2X1_7072 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10467) );
	NAND2X1 NAND2X1_7073 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10466), .B(dp.rf._abc_6362_n10467), .Y(dp.rf._abc_6362_n10468) );
	NAND2X1 NAND2X1_7074 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10468), .Y(dp.rf._abc_6362_n10469) );
	NAND2X1 NAND2X1_7075 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<20>), .Y(dp.rf._abc_6362_n10470) );
	NAND2X1 NAND2X1_7076 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10471) );
	NAND2X1 NAND2X1_7077 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10470), .B(dp.rf._abc_6362_n10471), .Y(dp.rf._abc_6362_n10472) );
	NAND2X1 NAND2X1_7078 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10472), .Y(dp.rf._abc_6362_n10473) );
	AND2X2 AND2X2_517 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10469), .B(dp.rf._abc_6362_n10473), .Y(dp.rf._abc_6362_n10474) );
	NAND2X1 NAND2X1_7079 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10474), .Y(dp.rf._abc_6362_n10475) );
	NAND2X1 NAND2X1_7080 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10475), .Y(dp.rf._abc_6362_n10476) );
	NOR2X1 NOR2X1_1314 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10465), .B(dp.rf._abc_6362_n10476), .Y(dp.rf._abc_6362_n10477) );
	NAND2X1 NAND2X1_7081 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<20>), .Y(dp.rf._abc_6362_n10478) );
	NAND2X1 NAND2X1_7082 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10478), .Y(dp.rf._abc_6362_n10479) );
	NOR2X1 NOR2X1_1315 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7390), .Y(dp.rf._abc_6362_n10480) );
	NOR2X1 NOR2X1_1316 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10479), .B(dp.rf._abc_6362_n10480), .Y(dp.rf._abc_6362_n10481) );
	NAND2X1 NAND2X1_7083 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<20>), .Y(dp.rf._abc_6362_n10482) );
	NAND2X1 NAND2X1_7084 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10482), .Y(dp.rf._abc_6362_n10483) );
	NOR2X1 NOR2X1_1317 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7395), .Y(dp.rf._abc_6362_n10484) );
	NOR2X1 NOR2X1_1318 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10483), .B(dp.rf._abc_6362_n10484), .Y(dp.rf._abc_6362_n10485) );
	OR2X2 OR2X2_112 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10481), .B(dp.rf._abc_6362_n10485), .Y(dp.rf._abc_6362_n10486) );
	NAND2X1 NAND2X1_7085 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10486), .Y(dp.rf._abc_6362_n10487) );
	NAND2X1 NAND2X1_7086 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<20>), .Y(dp.rf._abc_6362_n10488) );
	NAND2X1 NAND2X1_7087 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10488), .Y(dp.rf._abc_6362_n10489) );
	NOR2X1 NOR2X1_1319 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7402), .Y(dp.rf._abc_6362_n10490) );
	NOR2X1 NOR2X1_1320 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10489), .B(dp.rf._abc_6362_n10490), .Y(dp.rf._abc_6362_n10491) );
	NAND2X1 NAND2X1_7088 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<20>), .Y(dp.rf._abc_6362_n10492) );
	NAND2X1 NAND2X1_7089 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10492), .Y(dp.rf._abc_6362_n10493) );
	NOR2X1 NOR2X1_1321 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7407), .Y(dp.rf._abc_6362_n10494) );
	NOR2X1 NOR2X1_1322 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10493), .B(dp.rf._abc_6362_n10494), .Y(dp.rf._abc_6362_n10495) );
	OR2X2 OR2X2_113 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10491), .B(dp.rf._abc_6362_n10495), .Y(dp.rf._abc_6362_n10496) );
	NAND2X1 NAND2X1_7090 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10496), .Y(dp.rf._abc_6362_n10497) );
	AND2X2 AND2X2_518 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10497), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10498) );
	NAND2X1 NAND2X1_7091 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10487), .B(dp.rf._abc_6362_n10498), .Y(dp.rf._abc_6362_n10499) );
	NAND2X1 NAND2X1_7092 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10499), .Y(dp.rf._abc_6362_n10500) );
	NOR2X1 NOR2X1_1323 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10477), .B(dp.rf._abc_6362_n10500), .Y(dp.rf._abc_6362_n10501) );
	NAND2X1 NAND2X1_7093 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<20>), .Y(dp.rf._abc_6362_n10502) );
	NAND2X1 NAND2X1_7094 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10503) );
	NAND2X1 NAND2X1_7095 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10502), .B(dp.rf._abc_6362_n10503), .Y(dp.rf._abc_6362_n10504) );
	NAND2X1 NAND2X1_7096 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10504), .Y(dp.rf._abc_6362_n10505) );
	NAND2X1 NAND2X1_7097 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<20>), .Y(dp.rf._abc_6362_n10506) );
	NAND2X1 NAND2X1_7098 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10507) );
	NAND2X1 NAND2X1_7099 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10506), .B(dp.rf._abc_6362_n10507), .Y(dp.rf._abc_6362_n10508) );
	NAND2X1 NAND2X1_7100 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10508), .Y(dp.rf._abc_6362_n10509) );
	AND2X2 AND2X2_519 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10505), .B(dp.rf._abc_6362_n10509), .Y(dp.rf._abc_6362_n10510) );
	NAND2X1 NAND2X1_7101 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10510), .Y(dp.rf._abc_6362_n10511) );
	NAND2X1 NAND2X1_7102 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<20>), .Y(dp.rf._abc_6362_n10512) );
	NAND2X1 NAND2X1_7103 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10513) );
	NAND2X1 NAND2X1_7104 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10512), .B(dp.rf._abc_6362_n10513), .Y(dp.rf._abc_6362_n10514) );
	NAND2X1 NAND2X1_7105 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10514), .Y(dp.rf._abc_6362_n10515) );
	NAND2X1 NAND2X1_7106 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<20>), .Y(dp.rf._abc_6362_n10516) );
	NAND2X1 NAND2X1_7107 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10517) );
	NAND2X1 NAND2X1_7108 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10516), .B(dp.rf._abc_6362_n10517), .Y(dp.rf._abc_6362_n10518) );
	NAND2X1 NAND2X1_7109 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10518), .Y(dp.rf._abc_6362_n10519) );
	AND2X2 AND2X2_520 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10515), .B(dp.rf._abc_6362_n10519), .Y(dp.rf._abc_6362_n10520) );
	NAND2X1 NAND2X1_7110 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10520), .Y(dp.rf._abc_6362_n10521) );
	AND2X2 AND2X2_521 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10521), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10522) );
	NAND2X1 NAND2X1_7111 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10511), .B(dp.rf._abc_6362_n10522), .Y(dp.rf._abc_6362_n10523) );
	NAND2X1 NAND2X1_7112 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10524) );
	NAND2X1 NAND2X1_7113 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<20>), .Y(dp.rf._abc_6362_n10525) );
	AND2X2 AND2X2_522 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10525), .B(instr[17]), .Y(dp.rf._abc_6362_n10526) );
	NAND2X1 NAND2X1_7114 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10524), .B(dp.rf._abc_6362_n10526), .Y(dp.rf._abc_6362_n10527) );
	NAND2X1 NAND2X1_7115 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10528) );
	NAND2X1 NAND2X1_7116 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<20>), .Y(dp.rf._abc_6362_n10529) );
	AND2X2 AND2X2_523 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10529), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10530) );
	NAND2X1 NAND2X1_7117 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10528), .B(dp.rf._abc_6362_n10530), .Y(dp.rf._abc_6362_n10531) );
	NAND2X1 NAND2X1_7118 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10527), .B(dp.rf._abc_6362_n10531), .Y(dp.rf._abc_6362_n10532) );
	AND2X2 AND2X2_524 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10532), .B(instr[18]), .Y(dp.rf._abc_6362_n10533) );
	NAND2X1 NAND2X1_7119 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10534) );
	NAND2X1 NAND2X1_7120 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<20>), .Y(dp.rf._abc_6362_n10535) );
	AND2X2 AND2X2_525 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10535), .B(instr[17]), .Y(dp.rf._abc_6362_n10536) );
	NAND2X1 NAND2X1_7121 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10534), .B(dp.rf._abc_6362_n10536), .Y(dp.rf._abc_6362_n10537) );
	NAND2X1 NAND2X1_7122 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<20>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10538) );
	NAND2X1 NAND2X1_7123 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<20>), .Y(dp.rf._abc_6362_n10539) );
	AND2X2 AND2X2_526 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10539), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10540) );
	NAND2X1 NAND2X1_7124 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10538), .B(dp.rf._abc_6362_n10540), .Y(dp.rf._abc_6362_n10541) );
	NAND2X1 NAND2X1_7125 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10537), .B(dp.rf._abc_6362_n10541), .Y(dp.rf._abc_6362_n10542) );
	NAND2X1 NAND2X1_7126 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10542), .Y(dp.rf._abc_6362_n10543) );
	NAND2X1 NAND2X1_7127 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10543), .Y(dp.rf._abc_6362_n10544) );
	NOR2X1 NOR2X1_1324 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10533), .B(dp.rf._abc_6362_n10544), .Y(dp.rf._abc_6362_n10545) );
	NOR2X1 NOR2X1_1325 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10545), .Y(dp.rf._abc_6362_n10546) );
	NAND2X1 NAND2X1_7128 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10523), .B(dp.rf._abc_6362_n10546), .Y(dp.rf._abc_6362_n10547) );
	NAND2X1 NAND2X1_7129 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n10547), .Y(dp.rf._abc_6362_n10548) );
	NOR2X1 NOR2X1_1326 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10501), .B(dp.rf._abc_6362_n10548), .Y(writedata_20__RAW) );
	NAND2X1 NAND2X1_7130 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<21>), .Y(dp.rf._abc_6362_n10550) );
	NAND2X1 NAND2X1_7131 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10551) );
	NAND2X1 NAND2X1_7132 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10550), .B(dp.rf._abc_6362_n10551), .Y(dp.rf._abc_6362_n10552) );
	NAND2X1 NAND2X1_7133 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10552), .Y(dp.rf._abc_6362_n10553) );
	NAND2X1 NAND2X1_7134 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<21>), .Y(dp.rf._abc_6362_n10554) );
	NAND2X1 NAND2X1_7135 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10555) );
	NAND2X1 NAND2X1_7136 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10554), .B(dp.rf._abc_6362_n10555), .Y(dp.rf._abc_6362_n10556) );
	NAND2X1 NAND2X1_7137 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10556), .Y(dp.rf._abc_6362_n10557) );
	NAND2X1 NAND2X1_7138 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10553), .B(dp.rf._abc_6362_n10557), .Y(dp.rf._abc_6362_n10558) );
	NOR2X1 NOR2X1_1327 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10558), .Y(dp.rf._abc_6362_n10559) );
	NAND2X1 NAND2X1_7139 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<21>), .Y(dp.rf._abc_6362_n10560) );
	NAND2X1 NAND2X1_7140 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10561) );
	NAND2X1 NAND2X1_7141 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10560), .B(dp.rf._abc_6362_n10561), .Y(dp.rf._abc_6362_n10562) );
	NAND2X1 NAND2X1_7142 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10562), .Y(dp.rf._abc_6362_n10563) );
	NAND2X1 NAND2X1_7143 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<21>), .Y(dp.rf._abc_6362_n10564) );
	NAND2X1 NAND2X1_7144 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10565) );
	NAND2X1 NAND2X1_7145 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10564), .B(dp.rf._abc_6362_n10565), .Y(dp.rf._abc_6362_n10566) );
	NAND2X1 NAND2X1_7146 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10566), .Y(dp.rf._abc_6362_n10567) );
	AND2X2 AND2X2_527 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10563), .B(dp.rf._abc_6362_n10567), .Y(dp.rf._abc_6362_n10568) );
	NAND2X1 NAND2X1_7147 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10568), .Y(dp.rf._abc_6362_n10569) );
	NAND2X1 NAND2X1_7148 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n10569), .Y(dp.rf._abc_6362_n10570) );
	NOR2X1 NOR2X1_1328 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10559), .B(dp.rf._abc_6362_n10570), .Y(dp.rf._abc_6362_n10571) );
	NAND2X1 NAND2X1_7149 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<21>), .Y(dp.rf._abc_6362_n10572) );
	NAND2X1 NAND2X1_7150 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10573) );
	NAND2X1 NAND2X1_7151 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10572), .B(dp.rf._abc_6362_n10573), .Y(dp.rf._abc_6362_n10574) );
	NAND2X1 NAND2X1_7152 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10574), .Y(dp.rf._abc_6362_n10575) );
	NAND2X1 NAND2X1_7153 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<21>), .Y(dp.rf._abc_6362_n10576) );
	NAND2X1 NAND2X1_7154 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10577) );
	NAND2X1 NAND2X1_7155 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10576), .B(dp.rf._abc_6362_n10577), .Y(dp.rf._abc_6362_n10578) );
	NAND2X1 NAND2X1_7156 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10578), .Y(dp.rf._abc_6362_n10579) );
	NAND2X1 NAND2X1_7157 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10575), .B(dp.rf._abc_6362_n10579), .Y(dp.rf._abc_6362_n10580) );
	NAND2X1 NAND2X1_7158 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10580), .Y(dp.rf._abc_6362_n10581) );
	NAND2X1 NAND2X1_7159 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<21>), .Y(dp.rf._abc_6362_n10582) );
	NAND2X1 NAND2X1_7160 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10583) );
	NAND2X1 NAND2X1_7161 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10582), .B(dp.rf._abc_6362_n10583), .Y(dp.rf._abc_6362_n10584) );
	NAND2X1 NAND2X1_7162 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10584), .Y(dp.rf._abc_6362_n10585) );
	NAND2X1 NAND2X1_7163 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<21>), .Y(dp.rf._abc_6362_n10586) );
	NAND2X1 NAND2X1_7164 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10587) );
	NAND2X1 NAND2X1_7165 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10586), .B(dp.rf._abc_6362_n10587), .Y(dp.rf._abc_6362_n10588) );
	NAND2X1 NAND2X1_7166 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10588), .Y(dp.rf._abc_6362_n10589) );
	NAND2X1 NAND2X1_7167 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10585), .B(dp.rf._abc_6362_n10589), .Y(dp.rf._abc_6362_n10590) );
	NAND2X1 NAND2X1_7168 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10590), .Y(dp.rf._abc_6362_n10591) );
	NAND2X1 NAND2X1_7169 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10581), .B(dp.rf._abc_6362_n10591), .Y(dp.rf._abc_6362_n10592) );
	NAND2X1 NAND2X1_7170 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10592), .Y(dp.rf._abc_6362_n10593) );
	NAND2X1 NAND2X1_7171 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10593), .Y(dp.rf._abc_6362_n10594) );
	NOR2X1 NOR2X1_1329 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10571), .B(dp.rf._abc_6362_n10594), .Y(dp.rf._abc_6362_n10595) );
	NAND2X1 NAND2X1_7172 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<21>), .Y(dp.rf._abc_6362_n10596) );
	NAND2X1 NAND2X1_7173 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10596), .Y(dp.rf._abc_6362_n10597) );
	NOR2X1 NOR2X1_1330 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7513), .Y(dp.rf._abc_6362_n10598) );
	NOR2X1 NOR2X1_1331 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10597), .B(dp.rf._abc_6362_n10598), .Y(dp.rf._abc_6362_n10599) );
	NAND2X1 NAND2X1_7174 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<21>), .Y(dp.rf._abc_6362_n10600) );
	NAND2X1 NAND2X1_7175 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10600), .Y(dp.rf._abc_6362_n10601) );
	NOR2X1 NOR2X1_1332 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7518), .Y(dp.rf._abc_6362_n10602) );
	NOR2X1 NOR2X1_1333 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10601), .B(dp.rf._abc_6362_n10602), .Y(dp.rf._abc_6362_n10603) );
	OR2X2 OR2X2_114 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10599), .B(dp.rf._abc_6362_n10603), .Y(dp.rf._abc_6362_n10604) );
	NAND2X1 NAND2X1_7176 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10604), .Y(dp.rf._abc_6362_n10605) );
	NAND2X1 NAND2X1_7177 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<21>), .Y(dp.rf._abc_6362_n10606) );
	NAND2X1 NAND2X1_7178 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10606), .Y(dp.rf._abc_6362_n10607) );
	NOR2X1 NOR2X1_1334 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7525), .Y(dp.rf._abc_6362_n10608) );
	NOR2X1 NOR2X1_1335 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10607), .B(dp.rf._abc_6362_n10608), .Y(dp.rf._abc_6362_n10609) );
	NAND2X1 NAND2X1_7179 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<21>), .Y(dp.rf._abc_6362_n10610) );
	NAND2X1 NAND2X1_7180 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10610), .Y(dp.rf._abc_6362_n10611) );
	NOR2X1 NOR2X1_1336 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7530), .Y(dp.rf._abc_6362_n10612) );
	NOR2X1 NOR2X1_1337 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10611), .B(dp.rf._abc_6362_n10612), .Y(dp.rf._abc_6362_n10613) );
	OR2X2 OR2X2_115 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10609), .B(dp.rf._abc_6362_n10613), .Y(dp.rf._abc_6362_n10614) );
	NAND2X1 NAND2X1_7181 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10614), .Y(dp.rf._abc_6362_n10615) );
	AND2X2 AND2X2_528 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10615), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10616) );
	NAND2X1 NAND2X1_7182 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10605), .B(dp.rf._abc_6362_n10616), .Y(dp.rf._abc_6362_n10617) );
	NAND2X1 NAND2X1_7183 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10618) );
	NAND2X1 NAND2X1_7184 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<21>), .Y(dp.rf._abc_6362_n10619) );
	AND2X2 AND2X2_529 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10619), .B(instr[17]), .Y(dp.rf._abc_6362_n10620) );
	NAND2X1 NAND2X1_7185 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10618), .B(dp.rf._abc_6362_n10620), .Y(dp.rf._abc_6362_n10621) );
	NAND2X1 NAND2X1_7186 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10622) );
	NAND2X1 NAND2X1_7187 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<21>), .Y(dp.rf._abc_6362_n10623) );
	AND2X2 AND2X2_530 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10623), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10624) );
	NAND2X1 NAND2X1_7188 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10622), .B(dp.rf._abc_6362_n10624), .Y(dp.rf._abc_6362_n10625) );
	NAND2X1 NAND2X1_7189 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10621), .B(dp.rf._abc_6362_n10625), .Y(dp.rf._abc_6362_n10626) );
	AND2X2 AND2X2_531 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10626), .B(instr[18]), .Y(dp.rf._abc_6362_n10627) );
	NAND2X1 NAND2X1_7190 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10628) );
	NAND2X1 NAND2X1_7191 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<21>), .Y(dp.rf._abc_6362_n10629) );
	AND2X2 AND2X2_532 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10629), .B(instr[17]), .Y(dp.rf._abc_6362_n10630) );
	NAND2X1 NAND2X1_7192 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10628), .B(dp.rf._abc_6362_n10630), .Y(dp.rf._abc_6362_n10631) );
	NAND2X1 NAND2X1_7193 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<21>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10632) );
	NAND2X1 NAND2X1_7194 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<21>), .Y(dp.rf._abc_6362_n10633) );
	AND2X2 AND2X2_533 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10633), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10634) );
	NAND2X1 NAND2X1_7195 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10632), .B(dp.rf._abc_6362_n10634), .Y(dp.rf._abc_6362_n10635) );
	NAND2X1 NAND2X1_7196 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10631), .B(dp.rf._abc_6362_n10635), .Y(dp.rf._abc_6362_n10636) );
	NAND2X1 NAND2X1_7197 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10636), .Y(dp.rf._abc_6362_n10637) );
	NAND2X1 NAND2X1_7198 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10637), .Y(dp.rf._abc_6362_n10638) );
	NOR2X1 NOR2X1_1338 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10627), .B(dp.rf._abc_6362_n10638), .Y(dp.rf._abc_6362_n10639) );
	NOR2X1 NOR2X1_1339 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10639), .Y(dp.rf._abc_6362_n10640) );
	NAND2X1 NAND2X1_7199 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10617), .B(dp.rf._abc_6362_n10640), .Y(dp.rf._abc_6362_n10641) );
	NAND2X1 NAND2X1_7200 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n10641), .Y(dp.rf._abc_6362_n10642) );
	NOR2X1 NOR2X1_1340 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10595), .B(dp.rf._abc_6362_n10642), .Y(writedata_21__RAW) );
	NAND2X1 NAND2X1_7201 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<22>), .Y(dp.rf._abc_6362_n10644) );
	NAND2X1 NAND2X1_7202 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10644), .Y(dp.rf._abc_6362_n10645) );
	NOR2X1 NOR2X1_1341 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7565), .Y(dp.rf._abc_6362_n10646) );
	NOR2X1 NOR2X1_1342 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10645), .B(dp.rf._abc_6362_n10646), .Y(dp.rf._abc_6362_n10647) );
	NAND2X1 NAND2X1_7203 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<22>), .Y(dp.rf._abc_6362_n10648) );
	NAND2X1 NAND2X1_7204 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10648), .Y(dp.rf._abc_6362_n10649) );
	NOR2X1 NOR2X1_1343 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7570), .Y(dp.rf._abc_6362_n10650) );
	NOR2X1 NOR2X1_1344 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10649), .B(dp.rf._abc_6362_n10650), .Y(dp.rf._abc_6362_n10651) );
	NOR2X1 NOR2X1_1345 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10647), .B(dp.rf._abc_6362_n10651), .Y(dp.rf._abc_6362_n10652) );
	NAND2X1 NAND2X1_7205 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10652), .Y(dp.rf._abc_6362_n10653) );
	NAND2X1 NAND2X1_7206 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<22>), .Y(dp.rf._abc_6362_n10654) );
	NAND2X1 NAND2X1_7207 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10654), .Y(dp.rf._abc_6362_n10655) );
	NOR2X1 NOR2X1_1346 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7577), .Y(dp.rf._abc_6362_n10656) );
	NOR2X1 NOR2X1_1347 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10655), .B(dp.rf._abc_6362_n10656), .Y(dp.rf._abc_6362_n10657) );
	NAND2X1 NAND2X1_7208 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<22>), .Y(dp.rf._abc_6362_n10658) );
	NAND2X1 NAND2X1_7209 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10658), .Y(dp.rf._abc_6362_n10659) );
	NOR2X1 NOR2X1_1348 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7582), .Y(dp.rf._abc_6362_n10660) );
	NOR2X1 NOR2X1_1349 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10659), .B(dp.rf._abc_6362_n10660), .Y(dp.rf._abc_6362_n10661) );
	NOR2X1 NOR2X1_1350 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10657), .B(dp.rf._abc_6362_n10661), .Y(dp.rf._abc_6362_n10662) );
	NAND2X1 NAND2X1_7210 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10662), .Y(dp.rf._abc_6362_n10663) );
	NAND2X1 NAND2X1_7211 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10653), .B(dp.rf._abc_6362_n10663), .Y(dp.rf._abc_6362_n10664) );
	NAND2X1 NAND2X1_7212 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10664), .Y(dp.rf._abc_6362_n10665) );
	NAND2X1 NAND2X1_7213 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10665), .Y(dp.rf._abc_6362_n10666) );
	NAND2X1 NAND2X1_7214 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<22>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10667) );
	NOR2X1 NOR2X1_1351 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7591), .Y(dp.rf._abc_6362_n10668) );
	NOR2X1 NOR2X1_1352 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10668), .Y(dp.rf._abc_6362_n10669) );
	NAND2X1 NAND2X1_7215 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10667), .B(dp.rf._abc_6362_n10669), .Y(dp.rf._abc_6362_n10670) );
	NAND2X1 NAND2X1_7216 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<22>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10671) );
	NOR2X1 NOR2X1_1353 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7596), .Y(dp.rf._abc_6362_n10672) );
	NOR2X1 NOR2X1_1354 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10672), .Y(dp.rf._abc_6362_n10673) );
	NAND2X1 NAND2X1_7217 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10671), .B(dp.rf._abc_6362_n10673), .Y(dp.rf._abc_6362_n10674) );
	NAND2X1 NAND2X1_7218 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10670), .B(dp.rf._abc_6362_n10674), .Y(dp.rf._abc_6362_n10675) );
	NOR2X1 NOR2X1_1355 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10675), .Y(dp.rf._abc_6362_n10676) );
	NAND2X1 NAND2X1_7219 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<22>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10677) );
	NOR2X1 NOR2X1_1356 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7603), .Y(dp.rf._abc_6362_n10678) );
	NOR2X1 NOR2X1_1357 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10678), .Y(dp.rf._abc_6362_n10679) );
	NAND2X1 NAND2X1_7220 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10677), .B(dp.rf._abc_6362_n10679), .Y(dp.rf._abc_6362_n10680) );
	NAND2X1 NAND2X1_7221 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<22>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10681) );
	NOR2X1 NOR2X1_1358 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7608), .Y(dp.rf._abc_6362_n10682) );
	NOR2X1 NOR2X1_1359 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10682), .Y(dp.rf._abc_6362_n10683) );
	NAND2X1 NAND2X1_7222 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10681), .B(dp.rf._abc_6362_n10683), .Y(dp.rf._abc_6362_n10684) );
	NAND2X1 NAND2X1_7223 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10680), .B(dp.rf._abc_6362_n10684), .Y(dp.rf._abc_6362_n10685) );
	NOR2X1 NOR2X1_1360 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10685), .Y(dp.rf._abc_6362_n10686) );
	NOR2X1 NOR2X1_1361 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10676), .B(dp.rf._abc_6362_n10686), .Y(dp.rf._abc_6362_n10687) );
	NOR2X1 NOR2X1_1362 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10687), .Y(dp.rf._abc_6362_n10688) );
	NOR2X1 NOR2X1_1363 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10666), .B(dp.rf._abc_6362_n10688), .Y(dp.rf._abc_6362_n10689) );
	NAND2X1 NAND2X1_7224 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<22>), .Y(dp.rf._abc_6362_n10690) );
	NAND2X1 NAND2X1_7225 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10690), .Y(dp.rf._abc_6362_n10691) );
	NOR2X1 NOR2X1_1364 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7619), .Y(dp.rf._abc_6362_n10692) );
	NOR2X1 NOR2X1_1365 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10691), .B(dp.rf._abc_6362_n10692), .Y(dp.rf._abc_6362_n10693) );
	NAND2X1 NAND2X1_7226 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<22>), .Y(dp.rf._abc_6362_n10694) );
	NAND2X1 NAND2X1_7227 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10694), .Y(dp.rf._abc_6362_n10695) );
	NOR2X1 NOR2X1_1366 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7624), .Y(dp.rf._abc_6362_n10696) );
	NOR2X1 NOR2X1_1367 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10695), .B(dp.rf._abc_6362_n10696), .Y(dp.rf._abc_6362_n10697) );
	OR2X2 OR2X2_116 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10693), .B(dp.rf._abc_6362_n10697), .Y(dp.rf._abc_6362_n10698) );
	NAND2X1 NAND2X1_7228 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10698), .Y(dp.rf._abc_6362_n10699) );
	NAND2X1 NAND2X1_7229 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<22>), .Y(dp.rf._abc_6362_n10700) );
	NAND2X1 NAND2X1_7230 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10700), .Y(dp.rf._abc_6362_n10701) );
	NOR2X1 NOR2X1_1368 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7631), .Y(dp.rf._abc_6362_n10702) );
	NOR2X1 NOR2X1_1369 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10701), .B(dp.rf._abc_6362_n10702), .Y(dp.rf._abc_6362_n10703) );
	NAND2X1 NAND2X1_7231 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<22>), .Y(dp.rf._abc_6362_n10704) );
	NAND2X1 NAND2X1_7232 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10704), .Y(dp.rf._abc_6362_n10705) );
	NOR2X1 NOR2X1_1370 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7636), .Y(dp.rf._abc_6362_n10706) );
	NOR2X1 NOR2X1_1371 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10705), .B(dp.rf._abc_6362_n10706), .Y(dp.rf._abc_6362_n10707) );
	OR2X2 OR2X2_117 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10703), .B(dp.rf._abc_6362_n10707), .Y(dp.rf._abc_6362_n10708) );
	NAND2X1 NAND2X1_7233 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10708), .Y(dp.rf._abc_6362_n10709) );
	AND2X2 AND2X2_534 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10709), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10710) );
	NAND2X1 NAND2X1_7234 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10699), .B(dp.rf._abc_6362_n10710), .Y(dp.rf._abc_6362_n10711) );
	NAND2X1 NAND2X1_7235 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<22>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10712) );
	NAND2X1 NAND2X1_7236 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<22>), .Y(dp.rf._abc_6362_n10713) );
	AND2X2 AND2X2_535 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10713), .B(instr[17]), .Y(dp.rf._abc_6362_n10714) );
	NAND2X1 NAND2X1_7237 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10712), .B(dp.rf._abc_6362_n10714), .Y(dp.rf._abc_6362_n10715) );
	NAND2X1 NAND2X1_7238 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<22>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10716) );
	NAND2X1 NAND2X1_7239 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<22>), .Y(dp.rf._abc_6362_n10717) );
	AND2X2 AND2X2_536 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10717), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10718) );
	NAND2X1 NAND2X1_7240 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10716), .B(dp.rf._abc_6362_n10718), .Y(dp.rf._abc_6362_n10719) );
	NAND2X1 NAND2X1_7241 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10715), .B(dp.rf._abc_6362_n10719), .Y(dp.rf._abc_6362_n10720) );
	AND2X2 AND2X2_537 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10720), .B(instr[18]), .Y(dp.rf._abc_6362_n10721) );
	NAND2X1 NAND2X1_7242 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<22>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10722) );
	NAND2X1 NAND2X1_7243 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<22>), .Y(dp.rf._abc_6362_n10723) );
	AND2X2 AND2X2_538 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10723), .B(instr[17]), .Y(dp.rf._abc_6362_n10724) );
	NAND2X1 NAND2X1_7244 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10722), .B(dp.rf._abc_6362_n10724), .Y(dp.rf._abc_6362_n10725) );
	NAND2X1 NAND2X1_7245 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<22>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10726) );
	NAND2X1 NAND2X1_7246 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<22>), .Y(dp.rf._abc_6362_n10727) );
	AND2X2 AND2X2_539 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10727), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10728) );
	NAND2X1 NAND2X1_7247 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10726), .B(dp.rf._abc_6362_n10728), .Y(dp.rf._abc_6362_n10729) );
	NAND2X1 NAND2X1_7248 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10725), .B(dp.rf._abc_6362_n10729), .Y(dp.rf._abc_6362_n10730) );
	NAND2X1 NAND2X1_7249 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10730), .Y(dp.rf._abc_6362_n10731) );
	NAND2X1 NAND2X1_7250 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10731), .Y(dp.rf._abc_6362_n10732) );
	NOR2X1 NOR2X1_1372 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10721), .B(dp.rf._abc_6362_n10732), .Y(dp.rf._abc_6362_n10733) );
	NOR2X1 NOR2X1_1373 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10733), .Y(dp.rf._abc_6362_n10734) );
	NAND2X1 NAND2X1_7251 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10711), .B(dp.rf._abc_6362_n10734), .Y(dp.rf._abc_6362_n10735) );
	NAND2X1 NAND2X1_7252 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n10735), .Y(dp.rf._abc_6362_n10736) );
	NOR2X1 NOR2X1_1374 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10689), .B(dp.rf._abc_6362_n10736), .Y(writedata_22__RAW) );
	NAND2X1 NAND2X1_7253 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10738) );
	NOR2X1 NOR2X1_1375 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7697), .Y(dp.rf._abc_6362_n10739) );
	NOR2X1 NOR2X1_1376 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10739), .Y(dp.rf._abc_6362_n10740) );
	NAND2X1 NAND2X1_7254 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10738), .B(dp.rf._abc_6362_n10740), .Y(dp.rf._abc_6362_n10741) );
	NAND2X1 NAND2X1_7255 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10742) );
	NOR2X1 NOR2X1_1377 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7702), .Y(dp.rf._abc_6362_n10743) );
	NOR2X1 NOR2X1_1378 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10743), .Y(dp.rf._abc_6362_n10744) );
	NAND2X1 NAND2X1_7256 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10742), .B(dp.rf._abc_6362_n10744), .Y(dp.rf._abc_6362_n10745) );
	NAND2X1 NAND2X1_7257 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10741), .B(dp.rf._abc_6362_n10745), .Y(dp.rf._abc_6362_n10746) );
	NOR2X1 NOR2X1_1379 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10746), .Y(dp.rf._abc_6362_n10747) );
	NAND2X1 NAND2X1_7258 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10748) );
	NOR2X1 NOR2X1_1380 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7709), .Y(dp.rf._abc_6362_n10749) );
	NOR2X1 NOR2X1_1381 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10749), .Y(dp.rf._abc_6362_n10750) );
	NAND2X1 NAND2X1_7259 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10748), .B(dp.rf._abc_6362_n10750), .Y(dp.rf._abc_6362_n10751) );
	NAND2X1 NAND2X1_7260 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10752) );
	NOR2X1 NOR2X1_1382 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7714), .Y(dp.rf._abc_6362_n10753) );
	NOR2X1 NOR2X1_1383 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10753), .Y(dp.rf._abc_6362_n10754) );
	NAND2X1 NAND2X1_7261 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10752), .B(dp.rf._abc_6362_n10754), .Y(dp.rf._abc_6362_n10755) );
	NAND2X1 NAND2X1_7262 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10751), .B(dp.rf._abc_6362_n10755), .Y(dp.rf._abc_6362_n10756) );
	NOR2X1 NOR2X1_1384 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10756), .Y(dp.rf._abc_6362_n10757) );
	NOR2X1 NOR2X1_1385 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10747), .B(dp.rf._abc_6362_n10757), .Y(dp.rf._abc_6362_n10758) );
	NOR2X1 NOR2X1_1386 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10758), .Y(dp.rf._abc_6362_n10759) );
	NAND2X1 NAND2X1_7263 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<23>), .Y(dp.rf._abc_6362_n10760) );
	NAND2X1 NAND2X1_7264 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10760), .Y(dp.rf._abc_6362_n10761) );
	NOR2X1 NOR2X1_1387 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7683), .Y(dp.rf._abc_6362_n10762) );
	NOR2X1 NOR2X1_1388 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10761), .B(dp.rf._abc_6362_n10762), .Y(dp.rf._abc_6362_n10763) );
	NAND2X1 NAND2X1_7265 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<23>), .Y(dp.rf._abc_6362_n10764) );
	NAND2X1 NAND2X1_7266 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10764), .Y(dp.rf._abc_6362_n10765) );
	NOR2X1 NOR2X1_1389 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7688), .Y(dp.rf._abc_6362_n10766) );
	NOR2X1 NOR2X1_1390 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10765), .B(dp.rf._abc_6362_n10766), .Y(dp.rf._abc_6362_n10767) );
	OR2X2 OR2X2_118 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10763), .B(dp.rf._abc_6362_n10767), .Y(dp.rf._abc_6362_n10768) );
	NAND2X1 NAND2X1_7267 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10768), .Y(dp.rf._abc_6362_n10769) );
	NAND2X1 NAND2X1_7268 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<23>), .Y(dp.rf._abc_6362_n10770) );
	NAND2X1 NAND2X1_7269 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10770), .Y(dp.rf._abc_6362_n10771) );
	NOR2X1 NOR2X1_1391 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7671), .Y(dp.rf._abc_6362_n10772) );
	NOR2X1 NOR2X1_1392 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10771), .B(dp.rf._abc_6362_n10772), .Y(dp.rf._abc_6362_n10773) );
	NAND2X1 NAND2X1_7270 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<23>), .Y(dp.rf._abc_6362_n10774) );
	NAND2X1 NAND2X1_7271 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10774), .Y(dp.rf._abc_6362_n10775) );
	NOR2X1 NOR2X1_1393 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7676), .Y(dp.rf._abc_6362_n10776) );
	NOR2X1 NOR2X1_1394 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10775), .B(dp.rf._abc_6362_n10776), .Y(dp.rf._abc_6362_n10777) );
	OR2X2 OR2X2_119 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10773), .B(dp.rf._abc_6362_n10777), .Y(dp.rf._abc_6362_n10778) );
	NAND2X1 NAND2X1_7272 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10778), .Y(dp.rf._abc_6362_n10779) );
	AND2X2 AND2X2_540 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10779), .B(instr[19]), .Y(dp.rf._abc_6362_n10780) );
	NAND2X1 NAND2X1_7273 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10769), .B(dp.rf._abc_6362_n10780), .Y(dp.rf._abc_6362_n10781) );
	NAND2X1 NAND2X1_7274 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10781), .Y(dp.rf._abc_6362_n10782) );
	NOR2X1 NOR2X1_1395 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10759), .B(dp.rf._abc_6362_n10782), .Y(dp.rf._abc_6362_n10783) );
	NAND2X1 NAND2X1_7275 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<23>), .Y(dp.rf._abc_6362_n10784) );
	NAND2X1 NAND2X1_7276 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10785) );
	NAND2X1 NAND2X1_7277 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10784), .B(dp.rf._abc_6362_n10785), .Y(dp.rf._abc_6362_n10786) );
	NAND2X1 NAND2X1_7278 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10786), .Y(dp.rf._abc_6362_n10787) );
	NAND2X1 NAND2X1_7279 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<23>), .Y(dp.rf._abc_6362_n10788) );
	NAND2X1 NAND2X1_7280 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10789) );
	NAND2X1 NAND2X1_7281 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10788), .B(dp.rf._abc_6362_n10789), .Y(dp.rf._abc_6362_n10790) );
	NAND2X1 NAND2X1_7282 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10790), .Y(dp.rf._abc_6362_n10791) );
	NAND2X1 NAND2X1_7283 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10787), .B(dp.rf._abc_6362_n10791), .Y(dp.rf._abc_6362_n10792) );
	NAND2X1 NAND2X1_7284 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10792), .Y(dp.rf._abc_6362_n10793) );
	NAND2X1 NAND2X1_7285 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<23>), .Y(dp.rf._abc_6362_n10794) );
	NAND2X1 NAND2X1_7286 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10795) );
	NAND2X1 NAND2X1_7287 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10794), .B(dp.rf._abc_6362_n10795), .Y(dp.rf._abc_6362_n10796) );
	NAND2X1 NAND2X1_7288 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10796), .Y(dp.rf._abc_6362_n10797) );
	NAND2X1 NAND2X1_7289 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<23>), .Y(dp.rf._abc_6362_n10798) );
	NAND2X1 NAND2X1_7290 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10799) );
	NAND2X1 NAND2X1_7291 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10798), .B(dp.rf._abc_6362_n10799), .Y(dp.rf._abc_6362_n10800) );
	NAND2X1 NAND2X1_7292 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10800), .Y(dp.rf._abc_6362_n10801) );
	NAND2X1 NAND2X1_7293 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10797), .B(dp.rf._abc_6362_n10801), .Y(dp.rf._abc_6362_n10802) );
	NAND2X1 NAND2X1_7294 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10802), .Y(dp.rf._abc_6362_n10803) );
	NAND2X1 NAND2X1_7295 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10793), .B(dp.rf._abc_6362_n10803), .Y(dp.rf._abc_6362_n10804) );
	NAND2X1 NAND2X1_7296 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10804), .Y(dp.rf._abc_6362_n10805) );
	NAND2X1 NAND2X1_7297 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10806) );
	NAND2X1 NAND2X1_7298 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<23>), .Y(dp.rf._abc_6362_n10807) );
	AND2X2 AND2X2_541 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10807), .B(instr[17]), .Y(dp.rf._abc_6362_n10808) );
	NAND2X1 NAND2X1_7299 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10806), .B(dp.rf._abc_6362_n10808), .Y(dp.rf._abc_6362_n10809) );
	NAND2X1 NAND2X1_7300 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10810) );
	NAND2X1 NAND2X1_7301 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<23>), .Y(dp.rf._abc_6362_n10811) );
	AND2X2 AND2X2_542 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10811), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10812) );
	NAND2X1 NAND2X1_7302 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10810), .B(dp.rf._abc_6362_n10812), .Y(dp.rf._abc_6362_n10813) );
	NAND2X1 NAND2X1_7303 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10809), .B(dp.rf._abc_6362_n10813), .Y(dp.rf._abc_6362_n10814) );
	AND2X2 AND2X2_543 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10814), .B(instr[18]), .Y(dp.rf._abc_6362_n10815) );
	NAND2X1 NAND2X1_7304 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10816) );
	NAND2X1 NAND2X1_7305 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<23>), .Y(dp.rf._abc_6362_n10817) );
	AND2X2 AND2X2_544 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10817), .B(instr[17]), .Y(dp.rf._abc_6362_n10818) );
	NAND2X1 NAND2X1_7306 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10816), .B(dp.rf._abc_6362_n10818), .Y(dp.rf._abc_6362_n10819) );
	NAND2X1 NAND2X1_7307 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<23>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10820) );
	NAND2X1 NAND2X1_7308 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<23>), .Y(dp.rf._abc_6362_n10821) );
	AND2X2 AND2X2_545 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10821), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10822) );
	NAND2X1 NAND2X1_7309 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10820), .B(dp.rf._abc_6362_n10822), .Y(dp.rf._abc_6362_n10823) );
	NAND2X1 NAND2X1_7310 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10819), .B(dp.rf._abc_6362_n10823), .Y(dp.rf._abc_6362_n10824) );
	NAND2X1 NAND2X1_7311 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10824), .Y(dp.rf._abc_6362_n10825) );
	NAND2X1 NAND2X1_7312 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n10825), .Y(dp.rf._abc_6362_n10826) );
	NOR2X1 NOR2X1_1396 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10815), .B(dp.rf._abc_6362_n10826), .Y(dp.rf._abc_6362_n10827) );
	NOR2X1 NOR2X1_1397 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10827), .Y(dp.rf._abc_6362_n10828) );
	NAND2X1 NAND2X1_7313 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10805), .B(dp.rf._abc_6362_n10828), .Y(dp.rf._abc_6362_n10829) );
	NAND2X1 NAND2X1_7314 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n10829), .Y(dp.rf._abc_6362_n10830) );
	NOR2X1 NOR2X1_1398 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10783), .B(dp.rf._abc_6362_n10830), .Y(writedata_23__RAW) );
	NAND2X1 NAND2X1_7315 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10832) );
	NOR2X1 NOR2X1_1399 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7772), .Y(dp.rf._abc_6362_n10833) );
	NOR2X1 NOR2X1_1400 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10833), .Y(dp.rf._abc_6362_n10834) );
	NAND2X1 NAND2X1_7316 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10832), .B(dp.rf._abc_6362_n10834), .Y(dp.rf._abc_6362_n10835) );
	NAND2X1 NAND2X1_7317 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10836) );
	NOR2X1 NOR2X1_1401 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7777), .Y(dp.rf._abc_6362_n10837) );
	NOR2X1 NOR2X1_1402 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10837), .Y(dp.rf._abc_6362_n10838) );
	NAND2X1 NAND2X1_7318 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10836), .B(dp.rf._abc_6362_n10838), .Y(dp.rf._abc_6362_n10839) );
	NAND2X1 NAND2X1_7319 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10835), .B(dp.rf._abc_6362_n10839), .Y(dp.rf._abc_6362_n10840) );
	NAND2X1 NAND2X1_7320 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10840), .Y(dp.rf._abc_6362_n10841) );
	NAND2X1 NAND2X1_7321 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10842) );
	NOR2X1 NOR2X1_1403 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7784), .Y(dp.rf._abc_6362_n10843) );
	NOR2X1 NOR2X1_1404 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10843), .Y(dp.rf._abc_6362_n10844) );
	NAND2X1 NAND2X1_7322 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10842), .B(dp.rf._abc_6362_n10844), .Y(dp.rf._abc_6362_n10845) );
	NAND2X1 NAND2X1_7323 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10846) );
	NOR2X1 NOR2X1_1405 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7789), .Y(dp.rf._abc_6362_n10847) );
	NOR2X1 NOR2X1_1406 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10847), .Y(dp.rf._abc_6362_n10848) );
	NAND2X1 NAND2X1_7324 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10846), .B(dp.rf._abc_6362_n10848), .Y(dp.rf._abc_6362_n10849) );
	NAND2X1 NAND2X1_7325 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10845), .B(dp.rf._abc_6362_n10849), .Y(dp.rf._abc_6362_n10850) );
	NAND2X1 NAND2X1_7326 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10850), .Y(dp.rf._abc_6362_n10851) );
	NAND2X1 NAND2X1_7327 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10841), .B(dp.rf._abc_6362_n10851), .Y(dp.rf._abc_6362_n10852) );
	NOR2X1 NOR2X1_1407 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10852), .Y(dp.rf._abc_6362_n10853) );
	NAND2X1 NAND2X1_7328 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<24>), .Y(dp.rf._abc_6362_n10854) );
	NAND2X1 NAND2X1_7329 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10854), .Y(dp.rf._abc_6362_n10855) );
	NOR2X1 NOR2X1_1408 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7799), .Y(dp.rf._abc_6362_n10856) );
	NOR2X1 NOR2X1_1409 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10855), .B(dp.rf._abc_6362_n10856), .Y(dp.rf._abc_6362_n10857) );
	NAND2X1 NAND2X1_7330 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<24>), .Y(dp.rf._abc_6362_n10858) );
	NAND2X1 NAND2X1_7331 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10858), .Y(dp.rf._abc_6362_n10859) );
	NOR2X1 NOR2X1_1410 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7804), .Y(dp.rf._abc_6362_n10860) );
	NOR2X1 NOR2X1_1411 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10859), .B(dp.rf._abc_6362_n10860), .Y(dp.rf._abc_6362_n10861) );
	OR2X2 OR2X2_120 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10857), .B(dp.rf._abc_6362_n10861), .Y(dp.rf._abc_6362_n10862) );
	NAND2X1 NAND2X1_7332 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10862), .Y(dp.rf._abc_6362_n10863) );
	NAND2X1 NAND2X1_7333 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<24>), .Y(dp.rf._abc_6362_n10864) );
	NAND2X1 NAND2X1_7334 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10864), .Y(dp.rf._abc_6362_n10865) );
	NOR2X1 NOR2X1_1412 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7811), .Y(dp.rf._abc_6362_n10866) );
	NOR2X1 NOR2X1_1413 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10865), .B(dp.rf._abc_6362_n10866), .Y(dp.rf._abc_6362_n10867) );
	NAND2X1 NAND2X1_7335 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<24>), .Y(dp.rf._abc_6362_n10868) );
	NAND2X1 NAND2X1_7336 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10868), .Y(dp.rf._abc_6362_n10869) );
	NOR2X1 NOR2X1_1414 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7816), .Y(dp.rf._abc_6362_n10870) );
	NOR2X1 NOR2X1_1415 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10869), .B(dp.rf._abc_6362_n10870), .Y(dp.rf._abc_6362_n10871) );
	OR2X2 OR2X2_121 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10867), .B(dp.rf._abc_6362_n10871), .Y(dp.rf._abc_6362_n10872) );
	NAND2X1 NAND2X1_7337 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10872), .Y(dp.rf._abc_6362_n10873) );
	AND2X2 AND2X2_546 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10873), .B(instr[19]), .Y(dp.rf._abc_6362_n10874) );
	NAND2X1 NAND2X1_7338 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10863), .B(dp.rf._abc_6362_n10874), .Y(dp.rf._abc_6362_n10875) );
	NAND2X1 NAND2X1_7339 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10875), .Y(dp.rf._abc_6362_n10876) );
	NOR2X1 NOR2X1_1416 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10853), .B(dp.rf._abc_6362_n10876), .Y(dp.rf._abc_6362_n10877) );
	NAND2X1 NAND2X1_7340 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<24>), .Y(dp.rf._abc_6362_n10878) );
	NAND2X1 NAND2X1_7341 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10879) );
	NAND2X1 NAND2X1_7342 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10878), .B(dp.rf._abc_6362_n10879), .Y(dp.rf._abc_6362_n10880) );
	NAND2X1 NAND2X1_7343 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10880), .Y(dp.rf._abc_6362_n10881) );
	NAND2X1 NAND2X1_7344 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<24>), .Y(dp.rf._abc_6362_n10882) );
	NAND2X1 NAND2X1_7345 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10883) );
	NAND2X1 NAND2X1_7346 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10882), .B(dp.rf._abc_6362_n10883), .Y(dp.rf._abc_6362_n10884) );
	NAND2X1 NAND2X1_7347 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10884), .Y(dp.rf._abc_6362_n10885) );
	AND2X2 AND2X2_547 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10881), .B(dp.rf._abc_6362_n10885), .Y(dp.rf._abc_6362_n10886) );
	NAND2X1 NAND2X1_7348 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10886), .Y(dp.rf._abc_6362_n10887) );
	NAND2X1 NAND2X1_7349 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<24>), .Y(dp.rf._abc_6362_n10888) );
	NAND2X1 NAND2X1_7350 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10889) );
	NAND2X1 NAND2X1_7351 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10888), .B(dp.rf._abc_6362_n10889), .Y(dp.rf._abc_6362_n10890) );
	NAND2X1 NAND2X1_7352 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10890), .Y(dp.rf._abc_6362_n10891) );
	NAND2X1 NAND2X1_7353 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<24>), .Y(dp.rf._abc_6362_n10892) );
	NAND2X1 NAND2X1_7354 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10893) );
	NAND2X1 NAND2X1_7355 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10892), .B(dp.rf._abc_6362_n10893), .Y(dp.rf._abc_6362_n10894) );
	NAND2X1 NAND2X1_7356 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10894), .Y(dp.rf._abc_6362_n10895) );
	AND2X2 AND2X2_548 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10891), .B(dp.rf._abc_6362_n10895), .Y(dp.rf._abc_6362_n10896) );
	NAND2X1 NAND2X1_7357 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10896), .Y(dp.rf._abc_6362_n10897) );
	AND2X2 AND2X2_549 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10897), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n10898) );
	NAND2X1 NAND2X1_7358 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10887), .B(dp.rf._abc_6362_n10898), .Y(dp.rf._abc_6362_n10899) );
	NAND2X1 NAND2X1_7359 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10900) );
	NAND2X1 NAND2X1_7360 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<24>), .Y(dp.rf._abc_6362_n10901) );
	AND2X2 AND2X2_550 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10901), .B(instr[17]), .Y(dp.rf._abc_6362_n10902) );
	NAND2X1 NAND2X1_7361 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10900), .B(dp.rf._abc_6362_n10902), .Y(dp.rf._abc_6362_n10903) );
	NAND2X1 NAND2X1_7362 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10904) );
	NAND2X1 NAND2X1_7363 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<24>), .Y(dp.rf._abc_6362_n10905) );
	AND2X2 AND2X2_551 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10905), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10906) );
	NAND2X1 NAND2X1_7364 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10904), .B(dp.rf._abc_6362_n10906), .Y(dp.rf._abc_6362_n10907) );
	NAND2X1 NAND2X1_7365 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10903), .B(dp.rf._abc_6362_n10907), .Y(dp.rf._abc_6362_n10908) );
	AND2X2 AND2X2_552 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10908), .B(instr[18]), .Y(dp.rf._abc_6362_n10909) );
	NAND2X1 NAND2X1_7366 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10910) );
	NAND2X1 NAND2X1_7367 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<24>), .Y(dp.rf._abc_6362_n10911) );
	AND2X2 AND2X2_553 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10911), .B(instr[17]), .Y(dp.rf._abc_6362_n10912) );
	NAND2X1 NAND2X1_7368 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10910), .B(dp.rf._abc_6362_n10912), .Y(dp.rf._abc_6362_n10913) );
	NAND2X1 NAND2X1_7369 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<24>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10914) );
	NAND2X1 NAND2X1_7370 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<24>), .Y(dp.rf._abc_6362_n10915) );
	AND2X2 AND2X2_554 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10915), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n10916) );
	NAND2X1 NAND2X1_7371 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10914), .B(dp.rf._abc_6362_n10916), .Y(dp.rf._abc_6362_n10917) );
	NAND2X1 NAND2X1_7372 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10913), .B(dp.rf._abc_6362_n10917), .Y(dp.rf._abc_6362_n10918) );
	NAND2X1 NAND2X1_7373 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10918), .Y(dp.rf._abc_6362_n10919) );
	NAND2X1 NAND2X1_7374 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10919), .Y(dp.rf._abc_6362_n10920) );
	NOR2X1 NOR2X1_1417 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10909), .B(dp.rf._abc_6362_n10920), .Y(dp.rf._abc_6362_n10921) );
	NOR2X1 NOR2X1_1418 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10921), .Y(dp.rf._abc_6362_n10922) );
	NAND2X1 NAND2X1_7375 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10899), .B(dp.rf._abc_6362_n10922), .Y(dp.rf._abc_6362_n10923) );
	NAND2X1 NAND2X1_7376 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n10923), .Y(dp.rf._abc_6362_n10924) );
	NOR2X1 NOR2X1_1419 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10877), .B(dp.rf._abc_6362_n10924), .Y(writedata_24__RAW) );
	NAND2X1 NAND2X1_7377 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<25>), .Y(dp.rf._abc_6362_n10926) );
	NAND2X1 NAND2X1_7378 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10926), .Y(dp.rf._abc_6362_n10927) );
	NOR2X1 NOR2X1_1420 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7913), .Y(dp.rf._abc_6362_n10928) );
	NOR2X1 NOR2X1_1421 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10927), .B(dp.rf._abc_6362_n10928), .Y(dp.rf._abc_6362_n10929) );
	NAND2X1 NAND2X1_7379 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<25>), .Y(dp.rf._abc_6362_n10930) );
	NAND2X1 NAND2X1_7380 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10930), .Y(dp.rf._abc_6362_n10931) );
	NOR2X1 NOR2X1_1422 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7918), .Y(dp.rf._abc_6362_n10932) );
	NOR2X1 NOR2X1_1423 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10931), .B(dp.rf._abc_6362_n10932), .Y(dp.rf._abc_6362_n10933) );
	NOR2X1 NOR2X1_1424 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10929), .B(dp.rf._abc_6362_n10933), .Y(dp.rf._abc_6362_n10934) );
	NAND2X1 NAND2X1_7381 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10934), .Y(dp.rf._abc_6362_n10935) );
	NAND2X1 NAND2X1_7382 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<25>), .Y(dp.rf._abc_6362_n10936) );
	NAND2X1 NAND2X1_7383 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10936), .Y(dp.rf._abc_6362_n10937) );
	NOR2X1 NOR2X1_1425 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7901), .Y(dp.rf._abc_6362_n10938) );
	NOR2X1 NOR2X1_1426 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10937), .B(dp.rf._abc_6362_n10938), .Y(dp.rf._abc_6362_n10939) );
	NAND2X1 NAND2X1_7384 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<25>), .Y(dp.rf._abc_6362_n10940) );
	NAND2X1 NAND2X1_7385 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10940), .Y(dp.rf._abc_6362_n10941) );
	NOR2X1 NOR2X1_1427 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n7906), .Y(dp.rf._abc_6362_n10942) );
	NOR2X1 NOR2X1_1428 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10941), .B(dp.rf._abc_6362_n10942), .Y(dp.rf._abc_6362_n10943) );
	NOR2X1 NOR2X1_1429 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10939), .B(dp.rf._abc_6362_n10943), .Y(dp.rf._abc_6362_n10944) );
	NAND2X1 NAND2X1_7386 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10944), .Y(dp.rf._abc_6362_n10945) );
	NAND2X1 NAND2X1_7387 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10935), .B(dp.rf._abc_6362_n10945), .Y(dp.rf._abc_6362_n10946) );
	NAND2X1 NAND2X1_7388 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10946), .Y(dp.rf._abc_6362_n10947) );
	NAND2X1 NAND2X1_7389 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n10947), .Y(dp.rf._abc_6362_n10948) );
	NAND2X1 NAND2X1_7390 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10949) );
	NOR2X1 NOR2X1_1430 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7886), .Y(dp.rf._abc_6362_n10950) );
	NOR2X1 NOR2X1_1431 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10950), .Y(dp.rf._abc_6362_n10951) );
	NAND2X1 NAND2X1_7391 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10949), .B(dp.rf._abc_6362_n10951), .Y(dp.rf._abc_6362_n10952) );
	NAND2X1 NAND2X1_7392 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10953) );
	NOR2X1 NOR2X1_1432 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7891), .Y(dp.rf._abc_6362_n10954) );
	NOR2X1 NOR2X1_1433 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10954), .Y(dp.rf._abc_6362_n10955) );
	NAND2X1 NAND2X1_7393 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10953), .B(dp.rf._abc_6362_n10955), .Y(dp.rf._abc_6362_n10956) );
	NAND2X1 NAND2X1_7394 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10952), .B(dp.rf._abc_6362_n10956), .Y(dp.rf._abc_6362_n10957) );
	NOR2X1 NOR2X1_1434 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10957), .Y(dp.rf._abc_6362_n10958) );
	NAND2X1 NAND2X1_7395 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10959) );
	NOR2X1 NOR2X1_1435 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7874), .Y(dp.rf._abc_6362_n10960) );
	NOR2X1 NOR2X1_1436 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10960), .Y(dp.rf._abc_6362_n10961) );
	NAND2X1 NAND2X1_7396 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10959), .B(dp.rf._abc_6362_n10961), .Y(dp.rf._abc_6362_n10962) );
	NAND2X1 NAND2X1_7397 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10963) );
	NOR2X1 NOR2X1_1437 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf._abc_6362_n7879), .Y(dp.rf._abc_6362_n10964) );
	NOR2X1 NOR2X1_1438 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10964), .Y(dp.rf._abc_6362_n10965) );
	NAND2X1 NAND2X1_7398 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10963), .B(dp.rf._abc_6362_n10965), .Y(dp.rf._abc_6362_n10966) );
	NAND2X1 NAND2X1_7399 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10962), .B(dp.rf._abc_6362_n10966), .Y(dp.rf._abc_6362_n10967) );
	NOR2X1 NOR2X1_1439 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10967), .Y(dp.rf._abc_6362_n10968) );
	NOR2X1 NOR2X1_1440 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10958), .B(dp.rf._abc_6362_n10968), .Y(dp.rf._abc_6362_n10969) );
	NOR2X1 NOR2X1_1441 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n10969), .Y(dp.rf._abc_6362_n10970) );
	NOR2X1 NOR2X1_1442 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10948), .B(dp.rf._abc_6362_n10970), .Y(dp.rf._abc_6362_n10971) );
	NAND2X1 NAND2X1_7400 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<25>), .Y(dp.rf._abc_6362_n10972) );
	NAND2X1 NAND2X1_7401 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10973) );
	NAND2X1 NAND2X1_7402 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10972), .B(dp.rf._abc_6362_n10973), .Y(dp.rf._abc_6362_n10974) );
	NAND2X1 NAND2X1_7403 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10974), .Y(dp.rf._abc_6362_n10975) );
	NAND2X1 NAND2X1_7404 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<25>), .Y(dp.rf._abc_6362_n10976) );
	NAND2X1 NAND2X1_7405 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10977) );
	NAND2X1 NAND2X1_7406 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10976), .B(dp.rf._abc_6362_n10977), .Y(dp.rf._abc_6362_n10978) );
	NAND2X1 NAND2X1_7407 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10978), .Y(dp.rf._abc_6362_n10979) );
	AND2X2 AND2X2_555 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10975), .B(dp.rf._abc_6362_n10979), .Y(dp.rf._abc_6362_n10980) );
	NAND2X1 NAND2X1_7408 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n10980), .Y(dp.rf._abc_6362_n10981) );
	NAND2X1 NAND2X1_7409 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<25>), .Y(dp.rf._abc_6362_n10982) );
	NAND2X1 NAND2X1_7410 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10983) );
	NAND2X1 NAND2X1_7411 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10982), .B(dp.rf._abc_6362_n10983), .Y(dp.rf._abc_6362_n10984) );
	NAND2X1 NAND2X1_7412 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n10984), .Y(dp.rf._abc_6362_n10985) );
	NAND2X1 NAND2X1_7413 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<25>), .Y(dp.rf._abc_6362_n10986) );
	NAND2X1 NAND2X1_7414 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10987) );
	NAND2X1 NAND2X1_7415 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10986), .B(dp.rf._abc_6362_n10987), .Y(dp.rf._abc_6362_n10988) );
	NAND2X1 NAND2X1_7416 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n10988), .Y(dp.rf._abc_6362_n10989) );
	AND2X2 AND2X2_556 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10985), .B(dp.rf._abc_6362_n10989), .Y(dp.rf._abc_6362_n10990) );
	NAND2X1 NAND2X1_7417 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n10990), .Y(dp.rf._abc_6362_n10991) );
	AND2X2 AND2X2_557 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10991), .B(instr[19]), .Y(dp.rf._abc_6362_n10992) );
	NAND2X1 NAND2X1_7418 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10981), .B(dp.rf._abc_6362_n10992), .Y(dp.rf._abc_6362_n10993) );
	NAND2X1 NAND2X1_7419 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10994) );
	NAND2X1 NAND2X1_7420 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<25>), .Y(dp.rf._abc_6362_n10995) );
	AND2X2 AND2X2_558 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10995), .B(instr[17]), .Y(dp.rf._abc_6362_n10996) );
	NAND2X1 NAND2X1_7421 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10994), .B(dp.rf._abc_6362_n10996), .Y(dp.rf._abc_6362_n10997) );
	NAND2X1 NAND2X1_7422 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n10998) );
	NAND2X1 NAND2X1_7423 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<25>), .Y(dp.rf._abc_6362_n10999) );
	AND2X2 AND2X2_559 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10999), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11000) );
	NAND2X1 NAND2X1_7424 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10998), .B(dp.rf._abc_6362_n11000), .Y(dp.rf._abc_6362_n11001) );
	NAND2X1 NAND2X1_7425 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10997), .B(dp.rf._abc_6362_n11001), .Y(dp.rf._abc_6362_n11002) );
	AND2X2 AND2X2_560 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11002), .B(instr[18]), .Y(dp.rf._abc_6362_n11003) );
	NAND2X1 NAND2X1_7426 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11004) );
	NAND2X1 NAND2X1_7427 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<25>), .Y(dp.rf._abc_6362_n11005) );
	AND2X2 AND2X2_561 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11005), .B(instr[17]), .Y(dp.rf._abc_6362_n11006) );
	NAND2X1 NAND2X1_7428 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11004), .B(dp.rf._abc_6362_n11006), .Y(dp.rf._abc_6362_n11007) );
	NAND2X1 NAND2X1_7429 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<25>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11008) );
	NAND2X1 NAND2X1_7430 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<25>), .Y(dp.rf._abc_6362_n11009) );
	AND2X2 AND2X2_562 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11009), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11010) );
	NAND2X1 NAND2X1_7431 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11008), .B(dp.rf._abc_6362_n11010), .Y(dp.rf._abc_6362_n11011) );
	NAND2X1 NAND2X1_7432 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11007), .B(dp.rf._abc_6362_n11011), .Y(dp.rf._abc_6362_n11012) );
	NAND2X1 NAND2X1_7433 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11012), .Y(dp.rf._abc_6362_n11013) );
	NAND2X1 NAND2X1_7434 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n11013), .Y(dp.rf._abc_6362_n11014) );
	NOR2X1 NOR2X1_1443 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11003), .B(dp.rf._abc_6362_n11014), .Y(dp.rf._abc_6362_n11015) );
	NOR2X1 NOR2X1_1444 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11015), .Y(dp.rf._abc_6362_n11016) );
	NAND2X1 NAND2X1_7435 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10993), .B(dp.rf._abc_6362_n11016), .Y(dp.rf._abc_6362_n11017) );
	NAND2X1 NAND2X1_7436 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n11017), .Y(dp.rf._abc_6362_n11018) );
	NOR2X1 NOR2X1_1445 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n10971), .B(dp.rf._abc_6362_n11018), .Y(writedata_25__RAW) );
	NAND2X1 NAND2X1_7437 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<26>), .Y(dp.rf._abc_6362_n11020) );
	NAND2X1 NAND2X1_7438 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11021) );
	NAND2X1 NAND2X1_7439 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11020), .B(dp.rf._abc_6362_n11021), .Y(dp.rf._abc_6362_n11022) );
	NAND2X1 NAND2X1_7440 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11022), .Y(dp.rf._abc_6362_n11023) );
	NAND2X1 NAND2X1_7441 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<26>), .Y(dp.rf._abc_6362_n11024) );
	NAND2X1 NAND2X1_7442 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11025) );
	NAND2X1 NAND2X1_7443 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11024), .B(dp.rf._abc_6362_n11025), .Y(dp.rf._abc_6362_n11026) );
	NAND2X1 NAND2X1_7444 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11026), .Y(dp.rf._abc_6362_n11027) );
	NAND2X1 NAND2X1_7445 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11023), .B(dp.rf._abc_6362_n11027), .Y(dp.rf._abc_6362_n11028) );
	NOR2X1 NOR2X1_1446 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11028), .Y(dp.rf._abc_6362_n11029) );
	NAND2X1 NAND2X1_7446 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<26>), .Y(dp.rf._abc_6362_n11030) );
	NAND2X1 NAND2X1_7447 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11031) );
	NAND2X1 NAND2X1_7448 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11030), .B(dp.rf._abc_6362_n11031), .Y(dp.rf._abc_6362_n11032) );
	NAND2X1 NAND2X1_7449 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11032), .Y(dp.rf._abc_6362_n11033) );
	NAND2X1 NAND2X1_7450 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<26>), .Y(dp.rf._abc_6362_n11034) );
	NAND2X1 NAND2X1_7451 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11035) );
	NAND2X1 NAND2X1_7452 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11034), .B(dp.rf._abc_6362_n11035), .Y(dp.rf._abc_6362_n11036) );
	NAND2X1 NAND2X1_7453 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11036), .Y(dp.rf._abc_6362_n11037) );
	AND2X2 AND2X2_563 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11033), .B(dp.rf._abc_6362_n11037), .Y(dp.rf._abc_6362_n11038) );
	NAND2X1 NAND2X1_7454 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11038), .Y(dp.rf._abc_6362_n11039) );
	NAND2X1 NAND2X1_7455 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n11039), .Y(dp.rf._abc_6362_n11040) );
	NOR2X1 NOR2X1_1447 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11029), .B(dp.rf._abc_6362_n11040), .Y(dp.rf._abc_6362_n11041) );
	NAND2X1 NAND2X1_7456 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<26>), .Y(dp.rf._abc_6362_n11042) );
	NAND2X1 NAND2X1_7457 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11043) );
	NAND2X1 NAND2X1_7458 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11042), .B(dp.rf._abc_6362_n11043), .Y(dp.rf._abc_6362_n11044) );
	NAND2X1 NAND2X1_7459 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11044), .Y(dp.rf._abc_6362_n11045) );
	NAND2X1 NAND2X1_7460 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<26>), .Y(dp.rf._abc_6362_n11046) );
	NAND2X1 NAND2X1_7461 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11047) );
	NAND2X1 NAND2X1_7462 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11046), .B(dp.rf._abc_6362_n11047), .Y(dp.rf._abc_6362_n11048) );
	NAND2X1 NAND2X1_7463 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11048), .Y(dp.rf._abc_6362_n11049) );
	AND2X2 AND2X2_564 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11045), .B(dp.rf._abc_6362_n11049), .Y(dp.rf._abc_6362_n11050) );
	NAND2X1 NAND2X1_7464 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11050), .Y(dp.rf._abc_6362_n11051) );
	NAND2X1 NAND2X1_7465 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<26>), .Y(dp.rf._abc_6362_n11052) );
	NAND2X1 NAND2X1_7466 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11052), .Y(dp.rf._abc_6362_n11053) );
	AND2X2 AND2X2_565 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf.rf_2_<26>), .Y(dp.rf._abc_6362_n11054) );
	NOR2X1 NOR2X1_1448 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11053), .B(dp.rf._abc_6362_n11054), .Y(dp.rf._abc_6362_n11055) );
	NAND2X1 NAND2X1_7467 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<26>), .Y(dp.rf._abc_6362_n11056) );
	NAND2X1 NAND2X1_7468 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11056), .Y(dp.rf._abc_6362_n11057) );
	INVX1 INVX1_260 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<26>), .Y(dp.rf._abc_6362_n11058) );
	NOR2X1 NOR2X1_1449 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n11058), .Y(dp.rf._abc_6362_n11059) );
	NOR2X1 NOR2X1_1450 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11057), .B(dp.rf._abc_6362_n11059), .Y(dp.rf._abc_6362_n11060) );
	OR2X2 OR2X2_122 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11055), .B(dp.rf._abc_6362_n11060), .Y(dp.rf._abc_6362_n11061) );
	NAND2X1 NAND2X1_7469 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11061), .Y(dp.rf._abc_6362_n11062) );
	AND2X2 AND2X2_566 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11062), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n11063) );
	NAND2X1 NAND2X1_7470 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11051), .B(dp.rf._abc_6362_n11063), .Y(dp.rf._abc_6362_n11064) );
	NAND2X1 NAND2X1_7471 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11064), .Y(dp.rf._abc_6362_n11065) );
	NOR2X1 NOR2X1_1451 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11041), .B(dp.rf._abc_6362_n11065), .Y(dp.rf._abc_6362_n11066) );
	NAND2X1 NAND2X1_7472 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<26>), .Y(dp.rf._abc_6362_n11067) );
	NAND2X1 NAND2X1_7473 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11068) );
	NAND2X1 NAND2X1_7474 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11067), .B(dp.rf._abc_6362_n11068), .Y(dp.rf._abc_6362_n11069) );
	NAND2X1 NAND2X1_7475 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11069), .Y(dp.rf._abc_6362_n11070) );
	NAND2X1 NAND2X1_7476 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<26>), .Y(dp.rf._abc_6362_n11071) );
	NAND2X1 NAND2X1_7477 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11072) );
	NAND2X1 NAND2X1_7478 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11071), .B(dp.rf._abc_6362_n11072), .Y(dp.rf._abc_6362_n11073) );
	NAND2X1 NAND2X1_7479 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11073), .Y(dp.rf._abc_6362_n11074) );
	AND2X2 AND2X2_567 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11070), .B(dp.rf._abc_6362_n11074), .Y(dp.rf._abc_6362_n11075) );
	NAND2X1 NAND2X1_7480 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11075), .Y(dp.rf._abc_6362_n11076) );
	NAND2X1 NAND2X1_7481 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<26>), .Y(dp.rf._abc_6362_n11077) );
	NAND2X1 NAND2X1_7482 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11078) );
	NAND2X1 NAND2X1_7483 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11077), .B(dp.rf._abc_6362_n11078), .Y(dp.rf._abc_6362_n11079) );
	NAND2X1 NAND2X1_7484 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11079), .Y(dp.rf._abc_6362_n11080) );
	NAND2X1 NAND2X1_7485 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<26>), .Y(dp.rf._abc_6362_n11081) );
	NAND2X1 NAND2X1_7486 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11082) );
	NAND2X1 NAND2X1_7487 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11081), .B(dp.rf._abc_6362_n11082), .Y(dp.rf._abc_6362_n11083) );
	NAND2X1 NAND2X1_7488 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11083), .Y(dp.rf._abc_6362_n11084) );
	AND2X2 AND2X2_568 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11080), .B(dp.rf._abc_6362_n11084), .Y(dp.rf._abc_6362_n11085) );
	NAND2X1 NAND2X1_7489 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11085), .Y(dp.rf._abc_6362_n11086) );
	AND2X2 AND2X2_569 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11086), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n11087) );
	NAND2X1 NAND2X1_7490 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11076), .B(dp.rf._abc_6362_n11087), .Y(dp.rf._abc_6362_n11088) );
	NAND2X1 NAND2X1_7491 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11089) );
	NAND2X1 NAND2X1_7492 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<26>), .Y(dp.rf._abc_6362_n11090) );
	AND2X2 AND2X2_570 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11090), .B(instr[17]), .Y(dp.rf._abc_6362_n11091) );
	NAND2X1 NAND2X1_7493 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11089), .B(dp.rf._abc_6362_n11091), .Y(dp.rf._abc_6362_n11092) );
	NAND2X1 NAND2X1_7494 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11093) );
	NAND2X1 NAND2X1_7495 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<26>), .Y(dp.rf._abc_6362_n11094) );
	AND2X2 AND2X2_571 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11094), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11095) );
	NAND2X1 NAND2X1_7496 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11093), .B(dp.rf._abc_6362_n11095), .Y(dp.rf._abc_6362_n11096) );
	NAND2X1 NAND2X1_7497 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11092), .B(dp.rf._abc_6362_n11096), .Y(dp.rf._abc_6362_n11097) );
	AND2X2 AND2X2_572 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11097), .B(instr[18]), .Y(dp.rf._abc_6362_n11098) );
	NAND2X1 NAND2X1_7498 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11099) );
	NAND2X1 NAND2X1_7499 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<26>), .Y(dp.rf._abc_6362_n11100) );
	AND2X2 AND2X2_573 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11100), .B(instr[17]), .Y(dp.rf._abc_6362_n11101) );
	NAND2X1 NAND2X1_7500 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11099), .B(dp.rf._abc_6362_n11101), .Y(dp.rf._abc_6362_n11102) );
	NAND2X1 NAND2X1_7501 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<26>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11103) );
	NAND2X1 NAND2X1_7502 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<26>), .Y(dp.rf._abc_6362_n11104) );
	AND2X2 AND2X2_574 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11104), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11105) );
	NAND2X1 NAND2X1_7503 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11103), .B(dp.rf._abc_6362_n11105), .Y(dp.rf._abc_6362_n11106) );
	NAND2X1 NAND2X1_7504 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11102), .B(dp.rf._abc_6362_n11106), .Y(dp.rf._abc_6362_n11107) );
	NAND2X1 NAND2X1_7505 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11107), .Y(dp.rf._abc_6362_n11108) );
	NAND2X1 NAND2X1_7506 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n11108), .Y(dp.rf._abc_6362_n11109) );
	NOR2X1 NOR2X1_1452 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11098), .B(dp.rf._abc_6362_n11109), .Y(dp.rf._abc_6362_n11110) );
	NOR2X1 NOR2X1_1453 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11110), .Y(dp.rf._abc_6362_n11111) );
	NAND2X1 NAND2X1_7507 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11088), .B(dp.rf._abc_6362_n11111), .Y(dp.rf._abc_6362_n11112) );
	NAND2X1 NAND2X1_7508 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n11112), .Y(dp.rf._abc_6362_n11113) );
	NOR2X1 NOR2X1_1454 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11066), .B(dp.rf._abc_6362_n11113), .Y(writedata_26__RAW) );
	NAND2X1 NAND2X1_7509 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<27>), .Y(dp.rf._abc_6362_n11115) );
	NAND2X1 NAND2X1_7510 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<27>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11116) );
	NAND2X1 NAND2X1_7511 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11115), .B(dp.rf._abc_6362_n11116), .Y(dp.rf._abc_6362_n11117) );
	NAND2X1 NAND2X1_7512 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11117), .Y(dp.rf._abc_6362_n11118) );
	NAND2X1 NAND2X1_7513 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<27>), .Y(dp.rf._abc_6362_n11119) );
	NAND2X1 NAND2X1_7514 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<27>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11120) );
	NAND2X1 NAND2X1_7515 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11119), .B(dp.rf._abc_6362_n11120), .Y(dp.rf._abc_6362_n11121) );
	NAND2X1 NAND2X1_7516 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11121), .Y(dp.rf._abc_6362_n11122) );
	NAND2X1 NAND2X1_7517 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11118), .B(dp.rf._abc_6362_n11122), .Y(dp.rf._abc_6362_n11123) );
	NOR2X1 NOR2X1_1455 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11123), .Y(dp.rf._abc_6362_n11124) );
	NAND2X1 NAND2X1_7518 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<27>), .Y(dp.rf._abc_6362_n11125) );
	NAND2X1 NAND2X1_7519 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<27>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11126) );
	NAND2X1 NAND2X1_7520 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11125), .B(dp.rf._abc_6362_n11126), .Y(dp.rf._abc_6362_n11127) );
	NAND2X1 NAND2X1_7521 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11127), .Y(dp.rf._abc_6362_n11128) );
	NAND2X1 NAND2X1_7522 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<27>), .Y(dp.rf._abc_6362_n11129) );
	NAND2X1 NAND2X1_7523 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<27>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11130) );
	NAND2X1 NAND2X1_7524 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11129), .B(dp.rf._abc_6362_n11130), .Y(dp.rf._abc_6362_n11131) );
	NAND2X1 NAND2X1_7525 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11131), .Y(dp.rf._abc_6362_n11132) );
	AND2X2 AND2X2_575 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11128), .B(dp.rf._abc_6362_n11132), .Y(dp.rf._abc_6362_n11133) );
	NAND2X1 NAND2X1_7526 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11133), .Y(dp.rf._abc_6362_n11134) );
	NAND2X1 NAND2X1_7527 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n11134), .Y(dp.rf._abc_6362_n11135) );
	NOR2X1 NOR2X1_1456 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11124), .B(dp.rf._abc_6362_n11135), .Y(dp.rf._abc_6362_n11136) );
	NAND2X1 NAND2X1_7528 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<27>), .Y(dp.rf._abc_6362_n11137) );
	NAND2X1 NAND2X1_7529 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<27>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11138) );
	NAND2X1 NAND2X1_7530 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11137), .B(dp.rf._abc_6362_n11138), .Y(dp.rf._abc_6362_n11139) );
	NAND2X1 NAND2X1_7531 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11139), .Y(dp.rf._abc_6362_n11140) );
	NAND2X1 NAND2X1_7532 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<27>), .Y(dp.rf._abc_6362_n11141) );
	NAND2X1 NAND2X1_7533 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<27>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11142) );
	NAND2X1 NAND2X1_7534 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11141), .B(dp.rf._abc_6362_n11142), .Y(dp.rf._abc_6362_n11143) );
	NAND2X1 NAND2X1_7535 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11143), .Y(dp.rf._abc_6362_n11144) );
	AND2X2 AND2X2_576 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11140), .B(dp.rf._abc_6362_n11144), .Y(dp.rf._abc_6362_n11145) );
	NAND2X1 NAND2X1_7536 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11145), .Y(dp.rf._abc_6362_n11146) );
	NAND2X1 NAND2X1_7537 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<27>), .Y(dp.rf._abc_6362_n11147) );
	NAND2X1 NAND2X1_7538 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11147), .Y(dp.rf._abc_6362_n11148) );
	AND2X2 AND2X2_577 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf.rf_10_<27>), .Y(dp.rf._abc_6362_n11149) );
	NOR2X1 NOR2X1_1457 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11148), .B(dp.rf._abc_6362_n11149), .Y(dp.rf._abc_6362_n11150) );
	NAND2X1 NAND2X1_7539 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<27>), .Y(dp.rf._abc_6362_n11151) );
	NAND2X1 NAND2X1_7540 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11151), .Y(dp.rf._abc_6362_n11152) );
	INVX1 INVX1_261 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<27>), .Y(dp.rf._abc_6362_n11153) );
	NOR2X1 NOR2X1_1458 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n11153), .Y(dp.rf._abc_6362_n11154) );
	NOR2X1 NOR2X1_1459 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11152), .B(dp.rf._abc_6362_n11154), .Y(dp.rf._abc_6362_n11155) );
	OR2X2 OR2X2_123 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11150), .B(dp.rf._abc_6362_n11155), .Y(dp.rf._abc_6362_n11156) );
	NAND2X1 NAND2X1_7541 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11156), .Y(dp.rf._abc_6362_n11157) );
	AND2X2 AND2X2_578 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11157), .B(instr[19]), .Y(dp.rf._abc_6362_n11158) );
	NAND2X1 NAND2X1_7542 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11146), .B(dp.rf._abc_6362_n11158), .Y(dp.rf._abc_6362_n11159) );
	NAND2X1 NAND2X1_7543 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11159), .Y(dp.rf._abc_6362_n11160) );
	NOR2X1 NOR2X1_1460 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11136), .B(dp.rf._abc_6362_n11160), .Y(dp.rf._abc_6362_n11161) );
	NAND2X1 NAND2X1_7544 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<27>), .Y(dp.rf._abc_6362_n11162) );
	NAND2X1 NAND2X1_7545 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11162), .Y(dp.rf._abc_6362_n11163) );
	NOR2X1 NOR2X1_1461 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8118), .Y(dp.rf._abc_6362_n11164) );
	NOR2X1 NOR2X1_1462 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11163), .B(dp.rf._abc_6362_n11164), .Y(dp.rf._abc_6362_n11165) );
	NAND2X1 NAND2X1_7546 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<27>), .Y(dp.rf._abc_6362_n11166) );
	NAND2X1 NAND2X1_7547 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11166), .Y(dp.rf._abc_6362_n11167) );
	NOR2X1 NOR2X1_1463 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8123), .Y(dp.rf._abc_6362_n11168) );
	NOR2X1 NOR2X1_1464 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11167), .B(dp.rf._abc_6362_n11168), .Y(dp.rf._abc_6362_n11169) );
	OR2X2 OR2X2_124 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11165), .B(dp.rf._abc_6362_n11169), .Y(dp.rf._abc_6362_n11170) );
	NAND2X1 NAND2X1_7548 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11170), .Y(dp.rf._abc_6362_n11171) );
	NAND2X1 NAND2X1_7549 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<27>), .Y(dp.rf._abc_6362_n11172) );
	NAND2X1 NAND2X1_7550 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11172), .Y(dp.rf._abc_6362_n11173) );
	NOR2X1 NOR2X1_1465 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8130), .Y(dp.rf._abc_6362_n11174) );
	NOR2X1 NOR2X1_1466 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11173), .B(dp.rf._abc_6362_n11174), .Y(dp.rf._abc_6362_n11175) );
	NAND2X1 NAND2X1_7551 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<27>), .Y(dp.rf._abc_6362_n11176) );
	NAND2X1 NAND2X1_7552 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11176), .Y(dp.rf._abc_6362_n11177) );
	NOR2X1 NOR2X1_1467 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8135), .Y(dp.rf._abc_6362_n11178) );
	NOR2X1 NOR2X1_1468 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11177), .B(dp.rf._abc_6362_n11178), .Y(dp.rf._abc_6362_n11179) );
	OR2X2 OR2X2_125 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11175), .B(dp.rf._abc_6362_n11179), .Y(dp.rf._abc_6362_n11180) );
	NAND2X1 NAND2X1_7553 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11180), .Y(dp.rf._abc_6362_n11181) );
	AND2X2 AND2X2_579 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11181), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n11182) );
	NAND2X1 NAND2X1_7554 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11171), .B(dp.rf._abc_6362_n11182), .Y(dp.rf._abc_6362_n11183) );
	NAND2X1 NAND2X1_7555 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<27>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11184) );
	NAND2X1 NAND2X1_7556 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<27>), .Y(dp.rf._abc_6362_n11185) );
	AND2X2 AND2X2_580 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11185), .B(instr[17]), .Y(dp.rf._abc_6362_n11186) );
	NAND2X1 NAND2X1_7557 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11184), .B(dp.rf._abc_6362_n11186), .Y(dp.rf._abc_6362_n11187) );
	NAND2X1 NAND2X1_7558 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<27>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11188) );
	NAND2X1 NAND2X1_7559 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<27>), .Y(dp.rf._abc_6362_n11189) );
	AND2X2 AND2X2_581 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11189), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11190) );
	NAND2X1 NAND2X1_7560 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11188), .B(dp.rf._abc_6362_n11190), .Y(dp.rf._abc_6362_n11191) );
	NAND2X1 NAND2X1_7561 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11187), .B(dp.rf._abc_6362_n11191), .Y(dp.rf._abc_6362_n11192) );
	AND2X2 AND2X2_582 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11192), .B(instr[18]), .Y(dp.rf._abc_6362_n11193) );
	NAND2X1 NAND2X1_7562 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<27>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11194) );
	NAND2X1 NAND2X1_7563 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<27>), .Y(dp.rf._abc_6362_n11195) );
	AND2X2 AND2X2_583 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11195), .B(instr[17]), .Y(dp.rf._abc_6362_n11196) );
	NAND2X1 NAND2X1_7564 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11194), .B(dp.rf._abc_6362_n11196), .Y(dp.rf._abc_6362_n11197) );
	NAND2X1 NAND2X1_7565 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<27>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11198) );
	NAND2X1 NAND2X1_7566 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<27>), .Y(dp.rf._abc_6362_n11199) );
	AND2X2 AND2X2_584 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11199), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11200) );
	NAND2X1 NAND2X1_7567 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11198), .B(dp.rf._abc_6362_n11200), .Y(dp.rf._abc_6362_n11201) );
	NAND2X1 NAND2X1_7568 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11197), .B(dp.rf._abc_6362_n11201), .Y(dp.rf._abc_6362_n11202) );
	NAND2X1 NAND2X1_7569 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11202), .Y(dp.rf._abc_6362_n11203) );
	NAND2X1 NAND2X1_7570 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n11203), .Y(dp.rf._abc_6362_n11204) );
	NOR2X1 NOR2X1_1469 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11193), .B(dp.rf._abc_6362_n11204), .Y(dp.rf._abc_6362_n11205) );
	NOR2X1 NOR2X1_1470 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11205), .Y(dp.rf._abc_6362_n11206) );
	NAND2X1 NAND2X1_7571 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11183), .B(dp.rf._abc_6362_n11206), .Y(dp.rf._abc_6362_n11207) );
	NAND2X1 NAND2X1_7572 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n11207), .Y(dp.rf._abc_6362_n11208) );
	NOR2X1 NOR2X1_1471 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11161), .B(dp.rf._abc_6362_n11208), .Y(writedata_27__RAW) );
	NAND2X1 NAND2X1_7573 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<28>), .Y(dp.rf._abc_6362_n11210) );
	NAND2X1 NAND2X1_7574 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<28>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11211) );
	NAND2X1 NAND2X1_7575 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11210), .B(dp.rf._abc_6362_n11211), .Y(dp.rf._abc_6362_n11212) );
	NAND2X1 NAND2X1_7576 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11212), .Y(dp.rf._abc_6362_n11213) );
	NAND2X1 NAND2X1_7577 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<28>), .Y(dp.rf._abc_6362_n11214) );
	NAND2X1 NAND2X1_7578 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<28>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11215) );
	NAND2X1 NAND2X1_7579 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11214), .B(dp.rf._abc_6362_n11215), .Y(dp.rf._abc_6362_n11216) );
	NAND2X1 NAND2X1_7580 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11216), .Y(dp.rf._abc_6362_n11217) );
	NAND2X1 NAND2X1_7581 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11213), .B(dp.rf._abc_6362_n11217), .Y(dp.rf._abc_6362_n11218) );
	NOR2X1 NOR2X1_1472 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11218), .Y(dp.rf._abc_6362_n11219) );
	NAND2X1 NAND2X1_7582 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<28>), .Y(dp.rf._abc_6362_n11220) );
	NAND2X1 NAND2X1_7583 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<28>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11221) );
	NAND2X1 NAND2X1_7584 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11220), .B(dp.rf._abc_6362_n11221), .Y(dp.rf._abc_6362_n11222) );
	NAND2X1 NAND2X1_7585 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11222), .Y(dp.rf._abc_6362_n11223) );
	NAND2X1 NAND2X1_7586 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<28>), .Y(dp.rf._abc_6362_n11224) );
	NAND2X1 NAND2X1_7587 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<28>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11225) );
	NAND2X1 NAND2X1_7588 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11224), .B(dp.rf._abc_6362_n11225), .Y(dp.rf._abc_6362_n11226) );
	NAND2X1 NAND2X1_7589 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11226), .Y(dp.rf._abc_6362_n11227) );
	AND2X2 AND2X2_585 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11223), .B(dp.rf._abc_6362_n11227), .Y(dp.rf._abc_6362_n11228) );
	NAND2X1 NAND2X1_7590 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11228), .Y(dp.rf._abc_6362_n11229) );
	NAND2X1 NAND2X1_7591 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n11229), .Y(dp.rf._abc_6362_n11230) );
	NOR2X1 NOR2X1_1473 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11219), .B(dp.rf._abc_6362_n11230), .Y(dp.rf._abc_6362_n11231) );
	NAND2X1 NAND2X1_7592 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<28>), .Y(dp.rf._abc_6362_n11232) );
	NAND2X1 NAND2X1_7593 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<28>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11233) );
	NAND2X1 NAND2X1_7594 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11232), .B(dp.rf._abc_6362_n11233), .Y(dp.rf._abc_6362_n11234) );
	NAND2X1 NAND2X1_7595 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11234), .Y(dp.rf._abc_6362_n11235) );
	NAND2X1 NAND2X1_7596 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<28>), .Y(dp.rf._abc_6362_n11236) );
	NAND2X1 NAND2X1_7597 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<28>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11237) );
	NAND2X1 NAND2X1_7598 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11236), .B(dp.rf._abc_6362_n11237), .Y(dp.rf._abc_6362_n11238) );
	NAND2X1 NAND2X1_7599 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11238), .Y(dp.rf._abc_6362_n11239) );
	AND2X2 AND2X2_586 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11235), .B(dp.rf._abc_6362_n11239), .Y(dp.rf._abc_6362_n11240) );
	NAND2X1 NAND2X1_7600 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11240), .Y(dp.rf._abc_6362_n11241) );
	NAND2X1 NAND2X1_7601 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<28>), .Y(dp.rf._abc_6362_n11242) );
	NAND2X1 NAND2X1_7602 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11242), .Y(dp.rf._abc_6362_n11243) );
	AND2X2 AND2X2_587 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf.rf_2_<28>), .Y(dp.rf._abc_6362_n11244) );
	NOR2X1 NOR2X1_1474 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11243), .B(dp.rf._abc_6362_n11244), .Y(dp.rf._abc_6362_n11245) );
	NAND2X1 NAND2X1_7603 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<28>), .Y(dp.rf._abc_6362_n11246) );
	NAND2X1 NAND2X1_7604 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11246), .Y(dp.rf._abc_6362_n11247) );
	INVX1 INVX1_262 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<28>), .Y(dp.rf._abc_6362_n11248) );
	NOR2X1 NOR2X1_1475 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n11248), .Y(dp.rf._abc_6362_n11249) );
	NOR2X1 NOR2X1_1476 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11247), .B(dp.rf._abc_6362_n11249), .Y(dp.rf._abc_6362_n11250) );
	OR2X2 OR2X2_126 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11245), .B(dp.rf._abc_6362_n11250), .Y(dp.rf._abc_6362_n11251) );
	NAND2X1 NAND2X1_7605 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11251), .Y(dp.rf._abc_6362_n11252) );
	AND2X2 AND2X2_588 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11252), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n11253) );
	NAND2X1 NAND2X1_7606 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11241), .B(dp.rf._abc_6362_n11253), .Y(dp.rf._abc_6362_n11254) );
	NAND2X1 NAND2X1_7607 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11254), .Y(dp.rf._abc_6362_n11255) );
	NOR2X1 NOR2X1_1477 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11231), .B(dp.rf._abc_6362_n11255), .Y(dp.rf._abc_6362_n11256) );
	NAND2X1 NAND2X1_7608 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<28>), .Y(dp.rf._abc_6362_n11257) );
	NAND2X1 NAND2X1_7609 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11257), .Y(dp.rf._abc_6362_n11258) );
	NOR2X1 NOR2X1_1478 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8216), .Y(dp.rf._abc_6362_n11259) );
	NOR2X1 NOR2X1_1479 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11258), .B(dp.rf._abc_6362_n11259), .Y(dp.rf._abc_6362_n11260) );
	NAND2X1 NAND2X1_7610 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<28>), .Y(dp.rf._abc_6362_n11261) );
	NAND2X1 NAND2X1_7611 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11261), .Y(dp.rf._abc_6362_n11262) );
	NOR2X1 NOR2X1_1480 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8221), .Y(dp.rf._abc_6362_n11263) );
	NOR2X1 NOR2X1_1481 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11262), .B(dp.rf._abc_6362_n11263), .Y(dp.rf._abc_6362_n11264) );
	OR2X2 OR2X2_127 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11260), .B(dp.rf._abc_6362_n11264), .Y(dp.rf._abc_6362_n11265) );
	NAND2X1 NAND2X1_7612 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11265), .Y(dp.rf._abc_6362_n11266) );
	NAND2X1 NAND2X1_7613 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<28>), .Y(dp.rf._abc_6362_n11267) );
	NAND2X1 NAND2X1_7614 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11267), .Y(dp.rf._abc_6362_n11268) );
	NOR2X1 NOR2X1_1482 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8228), .Y(dp.rf._abc_6362_n11269) );
	NOR2X1 NOR2X1_1483 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11268), .B(dp.rf._abc_6362_n11269), .Y(dp.rf._abc_6362_n11270) );
	NAND2X1 NAND2X1_7615 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<28>), .Y(dp.rf._abc_6362_n11271) );
	NAND2X1 NAND2X1_7616 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11271), .Y(dp.rf._abc_6362_n11272) );
	NOR2X1 NOR2X1_1484 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8233), .Y(dp.rf._abc_6362_n11273) );
	NOR2X1 NOR2X1_1485 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11272), .B(dp.rf._abc_6362_n11273), .Y(dp.rf._abc_6362_n11274) );
	OR2X2 OR2X2_128 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11270), .B(dp.rf._abc_6362_n11274), .Y(dp.rf._abc_6362_n11275) );
	NAND2X1 NAND2X1_7617 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11275), .Y(dp.rf._abc_6362_n11276) );
	AND2X2 AND2X2_589 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11276), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n11277) );
	NAND2X1 NAND2X1_7618 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11266), .B(dp.rf._abc_6362_n11277), .Y(dp.rf._abc_6362_n11278) );
	NAND2X1 NAND2X1_7619 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<28>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11279) );
	NAND2X1 NAND2X1_7620 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<28>), .Y(dp.rf._abc_6362_n11280) );
	AND2X2 AND2X2_590 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11280), .B(instr[17]), .Y(dp.rf._abc_6362_n11281) );
	NAND2X1 NAND2X1_7621 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11279), .B(dp.rf._abc_6362_n11281), .Y(dp.rf._abc_6362_n11282) );
	NAND2X1 NAND2X1_7622 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<28>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11283) );
	NAND2X1 NAND2X1_7623 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<28>), .Y(dp.rf._abc_6362_n11284) );
	AND2X2 AND2X2_591 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11284), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11285) );
	NAND2X1 NAND2X1_7624 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11283), .B(dp.rf._abc_6362_n11285), .Y(dp.rf._abc_6362_n11286) );
	NAND2X1 NAND2X1_7625 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11282), .B(dp.rf._abc_6362_n11286), .Y(dp.rf._abc_6362_n11287) );
	AND2X2 AND2X2_592 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11287), .B(instr[18]), .Y(dp.rf._abc_6362_n11288) );
	NAND2X1 NAND2X1_7626 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<28>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11289) );
	NAND2X1 NAND2X1_7627 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<28>), .Y(dp.rf._abc_6362_n11290) );
	AND2X2 AND2X2_593 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11290), .B(instr[17]), .Y(dp.rf._abc_6362_n11291) );
	NAND2X1 NAND2X1_7628 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11289), .B(dp.rf._abc_6362_n11291), .Y(dp.rf._abc_6362_n11292) );
	NAND2X1 NAND2X1_7629 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<28>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11293) );
	NAND2X1 NAND2X1_7630 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<28>), .Y(dp.rf._abc_6362_n11294) );
	AND2X2 AND2X2_594 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11294), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11295) );
	NAND2X1 NAND2X1_7631 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11293), .B(dp.rf._abc_6362_n11295), .Y(dp.rf._abc_6362_n11296) );
	NAND2X1 NAND2X1_7632 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11292), .B(dp.rf._abc_6362_n11296), .Y(dp.rf._abc_6362_n11297) );
	NAND2X1 NAND2X1_7633 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11297), .Y(dp.rf._abc_6362_n11298) );
	NAND2X1 NAND2X1_7634 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n11298), .Y(dp.rf._abc_6362_n11299) );
	NOR2X1 NOR2X1_1486 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11288), .B(dp.rf._abc_6362_n11299), .Y(dp.rf._abc_6362_n11300) );
	NOR2X1 NOR2X1_1487 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11300), .Y(dp.rf._abc_6362_n11301) );
	NAND2X1 NAND2X1_7635 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11278), .B(dp.rf._abc_6362_n11301), .Y(dp.rf._abc_6362_n11302) );
	NAND2X1 NAND2X1_7636 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n11302), .Y(dp.rf._abc_6362_n11303) );
	NOR2X1 NOR2X1_1488 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11256), .B(dp.rf._abc_6362_n11303), .Y(writedata_28__RAW) );
	NAND2X1 NAND2X1_7637 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<29>), .Y(dp.rf._abc_6362_n11305) );
	NAND2X1 NAND2X1_7638 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11306) );
	NAND2X1 NAND2X1_7639 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11305), .B(dp.rf._abc_6362_n11306), .Y(dp.rf._abc_6362_n11307) );
	NAND2X1 NAND2X1_7640 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11307), .Y(dp.rf._abc_6362_n11308) );
	NAND2X1 NAND2X1_7641 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<29>), .Y(dp.rf._abc_6362_n11309) );
	NAND2X1 NAND2X1_7642 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11310) );
	NAND2X1 NAND2X1_7643 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11309), .B(dp.rf._abc_6362_n11310), .Y(dp.rf._abc_6362_n11311) );
	NAND2X1 NAND2X1_7644 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11311), .Y(dp.rf._abc_6362_n11312) );
	NAND2X1 NAND2X1_7645 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11308), .B(dp.rf._abc_6362_n11312), .Y(dp.rf._abc_6362_n11313) );
	NOR2X1 NOR2X1_1489 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11313), .Y(dp.rf._abc_6362_n11314) );
	NAND2X1 NAND2X1_7646 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<29>), .Y(dp.rf._abc_6362_n11315) );
	NAND2X1 NAND2X1_7647 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11316) );
	NAND2X1 NAND2X1_7648 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11315), .B(dp.rf._abc_6362_n11316), .Y(dp.rf._abc_6362_n11317) );
	NAND2X1 NAND2X1_7649 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11317), .Y(dp.rf._abc_6362_n11318) );
	NAND2X1 NAND2X1_7650 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<29>), .Y(dp.rf._abc_6362_n11319) );
	NAND2X1 NAND2X1_7651 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_2_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11320) );
	NAND2X1 NAND2X1_7652 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11319), .B(dp.rf._abc_6362_n11320), .Y(dp.rf._abc_6362_n11321) );
	NAND2X1 NAND2X1_7653 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11321), .Y(dp.rf._abc_6362_n11322) );
	AND2X2 AND2X2_595 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11318), .B(dp.rf._abc_6362_n11322), .Y(dp.rf._abc_6362_n11323) );
	NAND2X1 NAND2X1_7654 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11323), .Y(dp.rf._abc_6362_n11324) );
	NAND2X1 NAND2X1_7655 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n11324), .Y(dp.rf._abc_6362_n11325) );
	NOR2X1 NOR2X1_1490 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11314), .B(dp.rf._abc_6362_n11325), .Y(dp.rf._abc_6362_n11326) );
	NAND2X1 NAND2X1_7656 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<29>), .Y(dp.rf._abc_6362_n11327) );
	NAND2X1 NAND2X1_7657 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11328) );
	NAND2X1 NAND2X1_7658 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11327), .B(dp.rf._abc_6362_n11328), .Y(dp.rf._abc_6362_n11329) );
	NAND2X1 NAND2X1_7659 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11329), .Y(dp.rf._abc_6362_n11330) );
	NAND2X1 NAND2X1_7660 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<29>), .Y(dp.rf._abc_6362_n11331) );
	NAND2X1 NAND2X1_7661 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11332) );
	NAND2X1 NAND2X1_7662 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11331), .B(dp.rf._abc_6362_n11332), .Y(dp.rf._abc_6362_n11333) );
	NAND2X1 NAND2X1_7663 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11333), .Y(dp.rf._abc_6362_n11334) );
	NAND2X1 NAND2X1_7664 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11330), .B(dp.rf._abc_6362_n11334), .Y(dp.rf._abc_6362_n11335) );
	NAND2X1 NAND2X1_7665 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11335), .Y(dp.rf._abc_6362_n11336) );
	NAND2X1 NAND2X1_7666 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<29>), .Y(dp.rf._abc_6362_n11337) );
	NAND2X1 NAND2X1_7667 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11338) );
	NAND2X1 NAND2X1_7668 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11337), .B(dp.rf._abc_6362_n11338), .Y(dp.rf._abc_6362_n11339) );
	NAND2X1 NAND2X1_7669 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11339), .Y(dp.rf._abc_6362_n11340) );
	NAND2X1 NAND2X1_7670 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<29>), .Y(dp.rf._abc_6362_n11341) );
	NAND2X1 NAND2X1_7671 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11342) );
	NAND2X1 NAND2X1_7672 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11341), .B(dp.rf._abc_6362_n11342), .Y(dp.rf._abc_6362_n11343) );
	NAND2X1 NAND2X1_7673 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11343), .Y(dp.rf._abc_6362_n11344) );
	NAND2X1 NAND2X1_7674 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11340), .B(dp.rf._abc_6362_n11344), .Y(dp.rf._abc_6362_n11345) );
	NAND2X1 NAND2X1_7675 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11345), .Y(dp.rf._abc_6362_n11346) );
	NAND2X1 NAND2X1_7676 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11336), .B(dp.rf._abc_6362_n11346), .Y(dp.rf._abc_6362_n11347) );
	NAND2X1 NAND2X1_7677 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n11347), .Y(dp.rf._abc_6362_n11348) );
	NAND2X1 NAND2X1_7678 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11348), .Y(dp.rf._abc_6362_n11349) );
	NOR2X1 NOR2X1_1491 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11326), .B(dp.rf._abc_6362_n11349), .Y(dp.rf._abc_6362_n11350) );
	NAND2X1 NAND2X1_7679 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<29>), .Y(dp.rf._abc_6362_n11351) );
	NAND2X1 NAND2X1_7680 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11351), .Y(dp.rf._abc_6362_n11352) );
	NOR2X1 NOR2X1_1492 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8315), .Y(dp.rf._abc_6362_n11353) );
	NOR2X1 NOR2X1_1493 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11352), .B(dp.rf._abc_6362_n11353), .Y(dp.rf._abc_6362_n11354) );
	NAND2X1 NAND2X1_7681 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<29>), .Y(dp.rf._abc_6362_n11355) );
	NAND2X1 NAND2X1_7682 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11355), .Y(dp.rf._abc_6362_n11356) );
	NOR2X1 NOR2X1_1494 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8320), .Y(dp.rf._abc_6362_n11357) );
	NOR2X1 NOR2X1_1495 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11356), .B(dp.rf._abc_6362_n11357), .Y(dp.rf._abc_6362_n11358) );
	OR2X2 OR2X2_129 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11354), .B(dp.rf._abc_6362_n11358), .Y(dp.rf._abc_6362_n11359) );
	NAND2X1 NAND2X1_7683 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11359), .Y(dp.rf._abc_6362_n11360) );
	NAND2X1 NAND2X1_7684 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<29>), .Y(dp.rf._abc_6362_n11361) );
	NAND2X1 NAND2X1_7685 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11361), .Y(dp.rf._abc_6362_n11362) );
	NOR2X1 NOR2X1_1496 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8327), .Y(dp.rf._abc_6362_n11363) );
	NOR2X1 NOR2X1_1497 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11362), .B(dp.rf._abc_6362_n11363), .Y(dp.rf._abc_6362_n11364) );
	NAND2X1 NAND2X1_7686 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<29>), .Y(dp.rf._abc_6362_n11365) );
	NAND2X1 NAND2X1_7687 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11365), .Y(dp.rf._abc_6362_n11366) );
	NOR2X1 NOR2X1_1498 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8332), .Y(dp.rf._abc_6362_n11367) );
	NOR2X1 NOR2X1_1499 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11366), .B(dp.rf._abc_6362_n11367), .Y(dp.rf._abc_6362_n11368) );
	OR2X2 OR2X2_130 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11364), .B(dp.rf._abc_6362_n11368), .Y(dp.rf._abc_6362_n11369) );
	NAND2X1 NAND2X1_7688 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11369), .Y(dp.rf._abc_6362_n11370) );
	AND2X2 AND2X2_596 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11370), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n11371) );
	NAND2X1 NAND2X1_7689 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11360), .B(dp.rf._abc_6362_n11371), .Y(dp.rf._abc_6362_n11372) );
	NAND2X1 NAND2X1_7690 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11373) );
	NAND2X1 NAND2X1_7691 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<29>), .Y(dp.rf._abc_6362_n11374) );
	AND2X2 AND2X2_597 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11374), .B(instr[17]), .Y(dp.rf._abc_6362_n11375) );
	NAND2X1 NAND2X1_7692 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11373), .B(dp.rf._abc_6362_n11375), .Y(dp.rf._abc_6362_n11376) );
	NAND2X1 NAND2X1_7693 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11377) );
	NAND2X1 NAND2X1_7694 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<29>), .Y(dp.rf._abc_6362_n11378) );
	AND2X2 AND2X2_598 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11378), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11379) );
	NAND2X1 NAND2X1_7695 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11377), .B(dp.rf._abc_6362_n11379), .Y(dp.rf._abc_6362_n11380) );
	NAND2X1 NAND2X1_7696 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11376), .B(dp.rf._abc_6362_n11380), .Y(dp.rf._abc_6362_n11381) );
	AND2X2 AND2X2_599 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11381), .B(instr[18]), .Y(dp.rf._abc_6362_n11382) );
	NAND2X1 NAND2X1_7697 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11383) );
	NAND2X1 NAND2X1_7698 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<29>), .Y(dp.rf._abc_6362_n11384) );
	AND2X2 AND2X2_600 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11384), .B(instr[17]), .Y(dp.rf._abc_6362_n11385) );
	NAND2X1 NAND2X1_7699 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11383), .B(dp.rf._abc_6362_n11385), .Y(dp.rf._abc_6362_n11386) );
	NAND2X1 NAND2X1_7700 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<29>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11387) );
	NAND2X1 NAND2X1_7701 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<29>), .Y(dp.rf._abc_6362_n11388) );
	AND2X2 AND2X2_601 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11388), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11389) );
	NAND2X1 NAND2X1_7702 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11387), .B(dp.rf._abc_6362_n11389), .Y(dp.rf._abc_6362_n11390) );
	NAND2X1 NAND2X1_7703 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11386), .B(dp.rf._abc_6362_n11390), .Y(dp.rf._abc_6362_n11391) );
	NAND2X1 NAND2X1_7704 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11391), .Y(dp.rf._abc_6362_n11392) );
	NAND2X1 NAND2X1_7705 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n11392), .Y(dp.rf._abc_6362_n11393) );
	NOR2X1 NOR2X1_1500 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11382), .B(dp.rf._abc_6362_n11393), .Y(dp.rf._abc_6362_n11394) );
	NOR2X1 NOR2X1_1501 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11394), .Y(dp.rf._abc_6362_n11395) );
	NAND2X1 NAND2X1_7706 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11372), .B(dp.rf._abc_6362_n11395), .Y(dp.rf._abc_6362_n11396) );
	NAND2X1 NAND2X1_7707 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n11396), .Y(dp.rf._abc_6362_n11397) );
	NOR2X1 NOR2X1_1502 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11350), .B(dp.rf._abc_6362_n11397), .Y(writedata_29__RAW) );
	NAND2X1 NAND2X1_7708 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<30>), .Y(dp.rf._abc_6362_n11399) );
	NAND2X1 NAND2X1_7709 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_8_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11400) );
	NAND2X1 NAND2X1_7710 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11399), .B(dp.rf._abc_6362_n11400), .Y(dp.rf._abc_6362_n11401) );
	NAND2X1 NAND2X1_7711 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11401), .Y(dp.rf._abc_6362_n11402) );
	NAND2X1 NAND2X1_7712 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<30>), .Y(dp.rf._abc_6362_n11403) );
	NAND2X1 NAND2X1_7713 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_10_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11404) );
	NAND2X1 NAND2X1_7714 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11403), .B(dp.rf._abc_6362_n11404), .Y(dp.rf._abc_6362_n11405) );
	NAND2X1 NAND2X1_7715 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11405), .Y(dp.rf._abc_6362_n11406) );
	NAND2X1 NAND2X1_7716 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11402), .B(dp.rf._abc_6362_n11406), .Y(dp.rf._abc_6362_n11407) );
	NOR2X1 NOR2X1_1503 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11407), .Y(dp.rf._abc_6362_n11408) );
	NAND2X1 NAND2X1_7717 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<30>), .Y(dp.rf._abc_6362_n11409) );
	NAND2X1 NAND2X1_7718 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_12_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11410) );
	NAND2X1 NAND2X1_7719 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11409), .B(dp.rf._abc_6362_n11410), .Y(dp.rf._abc_6362_n11411) );
	NAND2X1 NAND2X1_7720 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11411), .Y(dp.rf._abc_6362_n11412) );
	NAND2X1 NAND2X1_7721 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<30>), .Y(dp.rf._abc_6362_n11413) );
	NAND2X1 NAND2X1_7722 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_14_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11414) );
	NAND2X1 NAND2X1_7723 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11413), .B(dp.rf._abc_6362_n11414), .Y(dp.rf._abc_6362_n11415) );
	NAND2X1 NAND2X1_7724 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11415), .Y(dp.rf._abc_6362_n11416) );
	AND2X2 AND2X2_602 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11412), .B(dp.rf._abc_6362_n11416), .Y(dp.rf._abc_6362_n11417) );
	NAND2X1 NAND2X1_7725 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11417), .Y(dp.rf._abc_6362_n11418) );
	NAND2X1 NAND2X1_7726 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n11418), .Y(dp.rf._abc_6362_n11419) );
	NOR2X1 NOR2X1_1504 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11408), .B(dp.rf._abc_6362_n11419), .Y(dp.rf._abc_6362_n11420) );
	NAND2X1 NAND2X1_7727 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<30>), .Y(dp.rf._abc_6362_n11421) );
	NAND2X1 NAND2X1_7728 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_4_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11422) );
	NAND2X1 NAND2X1_7729 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11421), .B(dp.rf._abc_6362_n11422), .Y(dp.rf._abc_6362_n11423) );
	NAND2X1 NAND2X1_7730 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11423), .Y(dp.rf._abc_6362_n11424) );
	NAND2X1 NAND2X1_7731 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<30>), .Y(dp.rf._abc_6362_n11425) );
	NAND2X1 NAND2X1_7732 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_6_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11426) );
	NAND2X1 NAND2X1_7733 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11425), .B(dp.rf._abc_6362_n11426), .Y(dp.rf._abc_6362_n11427) );
	NAND2X1 NAND2X1_7734 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11427), .Y(dp.rf._abc_6362_n11428) );
	AND2X2 AND2X2_603 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11424), .B(dp.rf._abc_6362_n11428), .Y(dp.rf._abc_6362_n11429) );
	NAND2X1 NAND2X1_7735 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11429), .Y(dp.rf._abc_6362_n11430) );
	NAND2X1 NAND2X1_7736 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<30>), .Y(dp.rf._abc_6362_n11431) );
	NAND2X1 NAND2X1_7737 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11431), .Y(dp.rf._abc_6362_n11432) );
	AND2X2 AND2X2_604 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8587), .B(dp.rf.rf_2_<30>), .Y(dp.rf._abc_6362_n11433) );
	NOR2X1 NOR2X1_1505 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11432), .B(dp.rf._abc_6362_n11433), .Y(dp.rf._abc_6362_n11434) );
	NAND2X1 NAND2X1_7738 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<30>), .Y(dp.rf._abc_6362_n11435) );
	NAND2X1 NAND2X1_7739 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11435), .Y(dp.rf._abc_6362_n11436) );
	INVX1 INVX1_263 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_0_<30>), .Y(dp.rf._abc_6362_n11437) );
	NOR2X1 NOR2X1_1506 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n11437), .Y(dp.rf._abc_6362_n11438) );
	NOR2X1 NOR2X1_1507 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11436), .B(dp.rf._abc_6362_n11438), .Y(dp.rf._abc_6362_n11439) );
	OR2X2 OR2X2_131 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11434), .B(dp.rf._abc_6362_n11439), .Y(dp.rf._abc_6362_n11440) );
	NAND2X1 NAND2X1_7740 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11440), .Y(dp.rf._abc_6362_n11441) );
	AND2X2 AND2X2_605 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11441), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n11442) );
	NAND2X1 NAND2X1_7741 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11430), .B(dp.rf._abc_6362_n11442), .Y(dp.rf._abc_6362_n11443) );
	NAND2X1 NAND2X1_7742 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11443), .Y(dp.rf._abc_6362_n11444) );
	NOR2X1 NOR2X1_1508 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11420), .B(dp.rf._abc_6362_n11444), .Y(dp.rf._abc_6362_n11445) );
	NAND2X1 NAND2X1_7743 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<30>), .Y(dp.rf._abc_6362_n11446) );
	NAND2X1 NAND2X1_7744 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11447) );
	NAND2X1 NAND2X1_7745 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11446), .B(dp.rf._abc_6362_n11447), .Y(dp.rf._abc_6362_n11448) );
	NAND2X1 NAND2X1_7746 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11448), .Y(dp.rf._abc_6362_n11449) );
	NAND2X1 NAND2X1_7747 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<30>), .Y(dp.rf._abc_6362_n11450) );
	NAND2X1 NAND2X1_7748 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11451) );
	NAND2X1 NAND2X1_7749 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11450), .B(dp.rf._abc_6362_n11451), .Y(dp.rf._abc_6362_n11452) );
	NAND2X1 NAND2X1_7750 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11452), .Y(dp.rf._abc_6362_n11453) );
	AND2X2 AND2X2_606 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11449), .B(dp.rf._abc_6362_n11453), .Y(dp.rf._abc_6362_n11454) );
	NAND2X1 NAND2X1_7751 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11454), .Y(dp.rf._abc_6362_n11455) );
	NAND2X1 NAND2X1_7752 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<30>), .Y(dp.rf._abc_6362_n11456) );
	NAND2X1 NAND2X1_7753 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11457) );
	NAND2X1 NAND2X1_7754 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11456), .B(dp.rf._abc_6362_n11457), .Y(dp.rf._abc_6362_n11458) );
	NAND2X1 NAND2X1_7755 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11458), .Y(dp.rf._abc_6362_n11459) );
	NAND2X1 NAND2X1_7756 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<30>), .Y(dp.rf._abc_6362_n11460) );
	NAND2X1 NAND2X1_7757 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11461) );
	NAND2X1 NAND2X1_7758 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11460), .B(dp.rf._abc_6362_n11461), .Y(dp.rf._abc_6362_n11462) );
	NAND2X1 NAND2X1_7759 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11462), .Y(dp.rf._abc_6362_n11463) );
	AND2X2 AND2X2_607 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11459), .B(dp.rf._abc_6362_n11463), .Y(dp.rf._abc_6362_n11464) );
	NAND2X1 NAND2X1_7760 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11464), .Y(dp.rf._abc_6362_n11465) );
	AND2X2 AND2X2_608 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11465), .B(instr[19]), .Y(dp.rf._abc_6362_n11466) );
	NAND2X1 NAND2X1_7761 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11455), .B(dp.rf._abc_6362_n11466), .Y(dp.rf._abc_6362_n11467) );
	NAND2X1 NAND2X1_7762 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11468) );
	NAND2X1 NAND2X1_7763 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<30>), .Y(dp.rf._abc_6362_n11469) );
	AND2X2 AND2X2_609 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11469), .B(instr[17]), .Y(dp.rf._abc_6362_n11470) );
	NAND2X1 NAND2X1_7764 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11468), .B(dp.rf._abc_6362_n11470), .Y(dp.rf._abc_6362_n11471) );
	NAND2X1 NAND2X1_7765 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11472) );
	NAND2X1 NAND2X1_7766 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<30>), .Y(dp.rf._abc_6362_n11473) );
	AND2X2 AND2X2_610 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11473), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11474) );
	NAND2X1 NAND2X1_7767 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11472), .B(dp.rf._abc_6362_n11474), .Y(dp.rf._abc_6362_n11475) );
	NAND2X1 NAND2X1_7768 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11471), .B(dp.rf._abc_6362_n11475), .Y(dp.rf._abc_6362_n11476) );
	AND2X2 AND2X2_611 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11476), .B(instr[18]), .Y(dp.rf._abc_6362_n11477) );
	NAND2X1 NAND2X1_7769 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11478) );
	NAND2X1 NAND2X1_7770 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<30>), .Y(dp.rf._abc_6362_n11479) );
	AND2X2 AND2X2_612 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11479), .B(instr[17]), .Y(dp.rf._abc_6362_n11480) );
	NAND2X1 NAND2X1_7771 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11478), .B(dp.rf._abc_6362_n11480), .Y(dp.rf._abc_6362_n11481) );
	NAND2X1 NAND2X1_7772 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<30>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11482) );
	NAND2X1 NAND2X1_7773 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<30>), .Y(dp.rf._abc_6362_n11483) );
	AND2X2 AND2X2_613 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11483), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11484) );
	NAND2X1 NAND2X1_7774 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11482), .B(dp.rf._abc_6362_n11484), .Y(dp.rf._abc_6362_n11485) );
	NAND2X1 NAND2X1_7775 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11481), .B(dp.rf._abc_6362_n11485), .Y(dp.rf._abc_6362_n11486) );
	NAND2X1 NAND2X1_7776 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11486), .Y(dp.rf._abc_6362_n11487) );
	NAND2X1 NAND2X1_7777 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8612), .B(dp.rf._abc_6362_n11487), .Y(dp.rf._abc_6362_n11488) );
	NOR2X1 NOR2X1_1509 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11477), .B(dp.rf._abc_6362_n11488), .Y(dp.rf._abc_6362_n11489) );
	NOR2X1 NOR2X1_1510 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11489), .Y(dp.rf._abc_6362_n11490) );
	NAND2X1 NAND2X1_7778 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11467), .B(dp.rf._abc_6362_n11490), .Y(dp.rf._abc_6362_n11491) );
	NAND2X1 NAND2X1_7779 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n11491), .Y(dp.rf._abc_6362_n11492) );
	NOR2X1 NOR2X1_1511 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11445), .B(dp.rf._abc_6362_n11492), .Y(writedata_30__RAW) );
	NAND2X1 NAND2X1_7780 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_11_<31>), .Y(dp.rf._abc_6362_n11494) );
	NAND2X1 NAND2X1_7781 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11494), .Y(dp.rf._abc_6362_n11495) );
	NOR2X1 NOR2X1_1512 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8461), .Y(dp.rf._abc_6362_n11496) );
	NOR2X1 NOR2X1_1513 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11495), .B(dp.rf._abc_6362_n11496), .Y(dp.rf._abc_6362_n11497) );
	NAND2X1 NAND2X1_7782 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_9_<31>), .Y(dp.rf._abc_6362_n11498) );
	NAND2X1 NAND2X1_7783 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11498), .Y(dp.rf._abc_6362_n11499) );
	NOR2X1 NOR2X1_1514 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8466), .Y(dp.rf._abc_6362_n11500) );
	NOR2X1 NOR2X1_1515 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11499), .B(dp.rf._abc_6362_n11500), .Y(dp.rf._abc_6362_n11501) );
	NOR2X1 NOR2X1_1516 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11497), .B(dp.rf._abc_6362_n11501), .Y(dp.rf._abc_6362_n11502) );
	NAND2X1 NAND2X1_7784 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11502), .Y(dp.rf._abc_6362_n11503) );
	NAND2X1 NAND2X1_7785 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_15_<31>), .Y(dp.rf._abc_6362_n11504) );
	NAND2X1 NAND2X1_7786 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11504), .Y(dp.rf._abc_6362_n11505) );
	NOR2X1 NOR2X1_1517 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8473), .Y(dp.rf._abc_6362_n11506) );
	NOR2X1 NOR2X1_1518 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11505), .B(dp.rf._abc_6362_n11506), .Y(dp.rf._abc_6362_n11507) );
	NAND2X1 NAND2X1_7787 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_13_<31>), .Y(dp.rf._abc_6362_n11508) );
	NAND2X1 NAND2X1_7788 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11508), .Y(dp.rf._abc_6362_n11509) );
	NOR2X1 NOR2X1_1519 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8478), .Y(dp.rf._abc_6362_n11510) );
	NOR2X1 NOR2X1_1520 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11509), .B(dp.rf._abc_6362_n11510), .Y(dp.rf._abc_6362_n11511) );
	NOR2X1 NOR2X1_1521 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11507), .B(dp.rf._abc_6362_n11511), .Y(dp.rf._abc_6362_n11512) );
	NAND2X1 NAND2X1_7789 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11512), .Y(dp.rf._abc_6362_n11513) );
	NAND2X1 NAND2X1_7790 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11503), .B(dp.rf._abc_6362_n11513), .Y(dp.rf._abc_6362_n11514) );
	NAND2X1 NAND2X1_7791 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n11514), .Y(dp.rf._abc_6362_n11515) );
	NAND2X1 NAND2X1_7792 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_7_<31>), .Y(dp.rf._abc_6362_n11516) );
	NAND2X1 NAND2X1_7793 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11516), .Y(dp.rf._abc_6362_n11517) );
	NOR2X1 NOR2X1_1522 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8487), .Y(dp.rf._abc_6362_n11518) );
	NOR2X1 NOR2X1_1523 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11517), .B(dp.rf._abc_6362_n11518), .Y(dp.rf._abc_6362_n11519) );
	NAND2X1 NAND2X1_7794 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_5_<31>), .Y(dp.rf._abc_6362_n11520) );
	NAND2X1 NAND2X1_7795 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11520), .Y(dp.rf._abc_6362_n11521) );
	NOR2X1 NOR2X1_1524 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8492), .Y(dp.rf._abc_6362_n11522) );
	NOR2X1 NOR2X1_1525 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11521), .B(dp.rf._abc_6362_n11522), .Y(dp.rf._abc_6362_n11523) );
	OR2X2 OR2X2_132 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11519), .B(dp.rf._abc_6362_n11523), .Y(dp.rf._abc_6362_n11524) );
	NAND2X1 NAND2X1_7796 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11524), .Y(dp.rf._abc_6362_n11525) );
	NAND2X1 NAND2X1_7797 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_3_<31>), .Y(dp.rf._abc_6362_n11526) );
	NAND2X1 NAND2X1_7798 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11526), .Y(dp.rf._abc_6362_n11527) );
	NOR2X1 NOR2X1_1526 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8499), .Y(dp.rf._abc_6362_n11528) );
	NOR2X1 NOR2X1_1527 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11527), .B(dp.rf._abc_6362_n11528), .Y(dp.rf._abc_6362_n11529) );
	NAND2X1 NAND2X1_7799 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_1_<31>), .Y(dp.rf._abc_6362_n11530) );
	NAND2X1 NAND2X1_7800 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11530), .Y(dp.rf._abc_6362_n11531) );
	NOR2X1 NOR2X1_1528 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf._abc_6362_n8504), .Y(dp.rf._abc_6362_n11532) );
	NOR2X1 NOR2X1_1529 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11531), .B(dp.rf._abc_6362_n11532), .Y(dp.rf._abc_6362_n11533) );
	OR2X2 OR2X2_133 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11529), .B(dp.rf._abc_6362_n11533), .Y(dp.rf._abc_6362_n11534) );
	NAND2X1 NAND2X1_7801 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11534), .Y(dp.rf._abc_6362_n11535) );
	AND2X2 AND2X2_614 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11535), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n11536) );
	NAND2X1 NAND2X1_7802 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11525), .B(dp.rf._abc_6362_n11536), .Y(dp.rf._abc_6362_n11537) );
	NAND2X1 NAND2X1_7803 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11515), .B(dp.rf._abc_6362_n11537), .Y(dp.rf._abc_6362_n11538) );
	NOR2X1 NOR2X1_1530 ( .gnd(gnd), .vdd(vdd), .A(instr[20]), .B(dp.rf._abc_6362_n11538), .Y(dp.rf._abc_6362_n11539) );
	NAND2X1 NAND2X1_7804 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_21_<31>), .Y(dp.rf._abc_6362_n11540) );
	NAND2X1 NAND2X1_7805 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_20_<31>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11541) );
	NAND2X1 NAND2X1_7806 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11540), .B(dp.rf._abc_6362_n11541), .Y(dp.rf._abc_6362_n11542) );
	NAND2X1 NAND2X1_7807 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11542), .Y(dp.rf._abc_6362_n11543) );
	NAND2X1 NAND2X1_7808 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_23_<31>), .Y(dp.rf._abc_6362_n11544) );
	NAND2X1 NAND2X1_7809 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_22_<31>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11545) );
	NAND2X1 NAND2X1_7810 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11544), .B(dp.rf._abc_6362_n11545), .Y(dp.rf._abc_6362_n11546) );
	NAND2X1 NAND2X1_7811 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11546), .Y(dp.rf._abc_6362_n11547) );
	AND2X2 AND2X2_615 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11543), .B(dp.rf._abc_6362_n11547), .Y(dp.rf._abc_6362_n11548) );
	NAND2X1 NAND2X1_7812 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.rf._abc_6362_n11548), .Y(dp.rf._abc_6362_n11549) );
	NAND2X1 NAND2X1_7813 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_17_<31>), .Y(dp.rf._abc_6362_n11550) );
	NAND2X1 NAND2X1_7814 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_16_<31>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11551) );
	NAND2X1 NAND2X1_7815 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11550), .B(dp.rf._abc_6362_n11551), .Y(dp.rf._abc_6362_n11552) );
	NAND2X1 NAND2X1_7816 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8567), .B(dp.rf._abc_6362_n11552), .Y(dp.rf._abc_6362_n11553) );
	NAND2X1 NAND2X1_7817 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_19_<31>), .Y(dp.rf._abc_6362_n11554) );
	NAND2X1 NAND2X1_7818 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_18_<31>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11555) );
	NAND2X1 NAND2X1_7819 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11554), .B(dp.rf._abc_6362_n11555), .Y(dp.rf._abc_6362_n11556) );
	NAND2X1 NAND2X1_7820 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.rf._abc_6362_n11556), .Y(dp.rf._abc_6362_n11557) );
	AND2X2 AND2X2_616 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11553), .B(dp.rf._abc_6362_n11557), .Y(dp.rf._abc_6362_n11558) );
	NAND2X1 NAND2X1_7821 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11558), .Y(dp.rf._abc_6362_n11559) );
	AND2X2 AND2X2_617 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11559), .B(dp.rf._abc_6362_n8612), .Y(dp.rf._abc_6362_n11560) );
	NAND2X1 NAND2X1_7822 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11549), .B(dp.rf._abc_6362_n11560), .Y(dp.rf._abc_6362_n11561) );
	NAND2X1 NAND2X1_7823 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_30_<31>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11562) );
	NAND2X1 NAND2X1_7824 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_31_<31>), .Y(dp.rf._abc_6362_n11563) );
	AND2X2 AND2X2_618 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11563), .B(instr[17]), .Y(dp.rf._abc_6362_n11564) );
	NAND2X1 NAND2X1_7825 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11562), .B(dp.rf._abc_6362_n11564), .Y(dp.rf._abc_6362_n11565) );
	NAND2X1 NAND2X1_7826 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_28_<31>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11566) );
	NAND2X1 NAND2X1_7827 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_29_<31>), .Y(dp.rf._abc_6362_n11567) );
	AND2X2 AND2X2_619 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11567), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11568) );
	NAND2X1 NAND2X1_7828 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11566), .B(dp.rf._abc_6362_n11568), .Y(dp.rf._abc_6362_n11569) );
	NAND2X1 NAND2X1_7829 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11565), .B(dp.rf._abc_6362_n11569), .Y(dp.rf._abc_6362_n11570) );
	AND2X2 AND2X2_620 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11570), .B(instr[18]), .Y(dp.rf._abc_6362_n11571) );
	NAND2X1 NAND2X1_7830 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_26_<31>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11572) );
	NAND2X1 NAND2X1_7831 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_27_<31>), .Y(dp.rf._abc_6362_n11573) );
	AND2X2 AND2X2_621 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11573), .B(instr[17]), .Y(dp.rf._abc_6362_n11574) );
	NAND2X1 NAND2X1_7832 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11572), .B(dp.rf._abc_6362_n11574), .Y(dp.rf._abc_6362_n11575) );
	NAND2X1 NAND2X1_7833 ( .gnd(gnd), .vdd(vdd), .A(dp.rf.rf_24_<31>), .B(dp.rf._abc_6362_n8587), .Y(dp.rf._abc_6362_n11576) );
	NAND2X1 NAND2X1_7834 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.rf.rf_25_<31>), .Y(dp.rf._abc_6362_n11577) );
	AND2X2 AND2X2_622 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11577), .B(dp.rf._abc_6362_n8567), .Y(dp.rf._abc_6362_n11578) );
	NAND2X1 NAND2X1_7835 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11576), .B(dp.rf._abc_6362_n11578), .Y(dp.rf._abc_6362_n11579) );
	NAND2X1 NAND2X1_7836 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11575), .B(dp.rf._abc_6362_n11579), .Y(dp.rf._abc_6362_n11580) );
	NAND2X1 NAND2X1_7837 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8562), .B(dp.rf._abc_6362_n11580), .Y(dp.rf._abc_6362_n11581) );
	NAND2X1 NAND2X1_7838 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.rf._abc_6362_n11581), .Y(dp.rf._abc_6362_n11582) );
	NOR2X1 NOR2X1_1531 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11571), .B(dp.rf._abc_6362_n11582), .Y(dp.rf._abc_6362_n11583) );
	NOR2X1 NOR2X1_1532 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8561), .B(dp.rf._abc_6362_n11583), .Y(dp.rf._abc_6362_n11584) );
	NAND2X1 NAND2X1_7839 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11561), .B(dp.rf._abc_6362_n11584), .Y(dp.rf._abc_6362_n11585) );
	NAND2X1 NAND2X1_7840 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n8615), .B(dp.rf._abc_6362_n11585), .Y(dp.rf._abc_6362_n11586) );
	NOR2X1 NOR2X1_1533 ( .gnd(gnd), .vdd(vdd), .A(dp.rf._abc_6362_n11539), .B(dp.rf._abc_6362_n11586), .Y(writedata_31__RAW) );
	DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3031), .Q(dp.rf.rf_0_<0>) );
	DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3033), .Q(dp.rf.rf_0_<1>) );
	DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3035), .Q(dp.rf.rf_0_<2>) );
	DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3037), .Q(dp.rf.rf_0_<3>) );
	DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3039), .Q(dp.rf.rf_0_<4>) );
	DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3041), .Q(dp.rf.rf_0_<5>) );
	DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3043), .Q(dp.rf.rf_0_<6>) );
	DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3045), .Q(dp.rf.rf_0_<7>) );
	DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3047), .Q(dp.rf.rf_0_<8>) );
	DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3049), .Q(dp.rf.rf_0_<9>) );
	DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3051), .Q(dp.rf.rf_0_<10>) );
	DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3053), .Q(dp.rf.rf_0_<11>) );
	DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3055), .Q(dp.rf.rf_0_<12>) );
	DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3057), .Q(dp.rf.rf_0_<13>) );
	DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3059), .Q(dp.rf.rf_0_<14>) );
	DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3061), .Q(dp.rf.rf_0_<15>) );
	DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3063), .Q(dp.rf.rf_0_<16>) );
	DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3065), .Q(dp.rf.rf_0_<17>) );
	DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3067), .Q(dp.rf.rf_0_<18>) );
	DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3069), .Q(dp.rf.rf_0_<19>) );
	DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3071), .Q(dp.rf.rf_0_<20>) );
	DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3073), .Q(dp.rf.rf_0_<21>) );
	DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3075), .Q(dp.rf.rf_0_<22>) );
	DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3077), .Q(dp.rf.rf_0_<23>) );
	DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3079), .Q(dp.rf.rf_0_<24>) );
	DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3081), .Q(dp.rf.rf_0_<25>) );
	DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3083), .Q(dp.rf.rf_0_<26>) );
	DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3085), .Q(dp.rf.rf_0_<27>) );
	DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3087), .Q(dp.rf.rf_0_<28>) );
	DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3089), .Q(dp.rf.rf_0_<29>) );
	DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3091), .Q(dp.rf.rf_0_<30>) );
	DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3093), .Q(dp.rf.rf_0_<31>) );
	DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3094), .Q(dp.rf.rf_10_<0>) );
	DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3095), .Q(dp.rf.rf_10_<1>) );
	DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3096), .Q(dp.rf.rf_10_<2>) );
	DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3097), .Q(dp.rf.rf_10_<3>) );
	DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3098), .Q(dp.rf.rf_10_<4>) );
	DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3099), .Q(dp.rf.rf_10_<5>) );
	DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3100), .Q(dp.rf.rf_10_<6>) );
	DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3101), .Q(dp.rf.rf_10_<7>) );
	DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3102), .Q(dp.rf.rf_10_<8>) );
	DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3103), .Q(dp.rf.rf_10_<9>) );
	DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3104), .Q(dp.rf.rf_10_<10>) );
	DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3105), .Q(dp.rf.rf_10_<11>) );
	DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3106), .Q(dp.rf.rf_10_<12>) );
	DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3107), .Q(dp.rf.rf_10_<13>) );
	DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3108), .Q(dp.rf.rf_10_<14>) );
	DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3109), .Q(dp.rf.rf_10_<15>) );
	DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3110), .Q(dp.rf.rf_10_<16>) );
	DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3111), .Q(dp.rf.rf_10_<17>) );
	DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3112), .Q(dp.rf.rf_10_<18>) );
	DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3113), .Q(dp.rf.rf_10_<19>) );
	DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3114), .Q(dp.rf.rf_10_<20>) );
	DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3115), .Q(dp.rf.rf_10_<21>) );
	DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3116), .Q(dp.rf.rf_10_<22>) );
	DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3117), .Q(dp.rf.rf_10_<23>) );
	DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3118), .Q(dp.rf.rf_10_<24>) );
	DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3119), .Q(dp.rf.rf_10_<25>) );
	DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3120), .Q(dp.rf.rf_10_<26>) );
	DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3121), .Q(dp.rf.rf_10_<27>) );
	DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3122), .Q(dp.rf.rf_10_<28>) );
	DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3123), .Q(dp.rf.rf_10_<29>) );
	DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3124), .Q(dp.rf.rf_10_<30>) );
	DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3125), .Q(dp.rf.rf_10_<31>) );
	DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3126), .Q(dp.rf.rf_11_<0>) );
	DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3127), .Q(dp.rf.rf_11_<1>) );
	DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3128), .Q(dp.rf.rf_11_<2>) );
	DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3129), .Q(dp.rf.rf_11_<3>) );
	DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3130), .Q(dp.rf.rf_11_<4>) );
	DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3131), .Q(dp.rf.rf_11_<5>) );
	DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3132), .Q(dp.rf.rf_11_<6>) );
	DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3133), .Q(dp.rf.rf_11_<7>) );
	DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3134), .Q(dp.rf.rf_11_<8>) );
	DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3135), .Q(dp.rf.rf_11_<9>) );
	DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3136), .Q(dp.rf.rf_11_<10>) );
	DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3137), .Q(dp.rf.rf_11_<11>) );
	DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3138), .Q(dp.rf.rf_11_<12>) );
	DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3139), .Q(dp.rf.rf_11_<13>) );
	DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3140), .Q(dp.rf.rf_11_<14>) );
	DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3141), .Q(dp.rf.rf_11_<15>) );
	DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3142), .Q(dp.rf.rf_11_<16>) );
	DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3143), .Q(dp.rf.rf_11_<17>) );
	DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3144), .Q(dp.rf.rf_11_<18>) );
	DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3145), .Q(dp.rf.rf_11_<19>) );
	DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3146), .Q(dp.rf.rf_11_<20>) );
	DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3147), .Q(dp.rf.rf_11_<21>) );
	DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3148), .Q(dp.rf.rf_11_<22>) );
	DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3149), .Q(dp.rf.rf_11_<23>) );
	DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3150), .Q(dp.rf.rf_11_<24>) );
	DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3151), .Q(dp.rf.rf_11_<25>) );
	DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3152), .Q(dp.rf.rf_11_<26>) );
	DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3153), .Q(dp.rf.rf_11_<27>) );
	DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3154), .Q(dp.rf.rf_11_<28>) );
	DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3155), .Q(dp.rf.rf_11_<29>) );
	DFFPOSX1 DFFPOSX1_95 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3156), .Q(dp.rf.rf_11_<30>) );
	DFFPOSX1 DFFPOSX1_96 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3157), .Q(dp.rf.rf_11_<31>) );
	DFFPOSX1 DFFPOSX1_97 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3158), .Q(dp.rf.rf_12_<0>) );
	DFFPOSX1 DFFPOSX1_98 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3159), .Q(dp.rf.rf_12_<1>) );
	DFFPOSX1 DFFPOSX1_99 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3160), .Q(dp.rf.rf_12_<2>) );
	DFFPOSX1 DFFPOSX1_100 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3161), .Q(dp.rf.rf_12_<3>) );
	DFFPOSX1 DFFPOSX1_101 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3162), .Q(dp.rf.rf_12_<4>) );
	DFFPOSX1 DFFPOSX1_102 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3163), .Q(dp.rf.rf_12_<5>) );
	DFFPOSX1 DFFPOSX1_103 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3164), .Q(dp.rf.rf_12_<6>) );
	DFFPOSX1 DFFPOSX1_104 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3165), .Q(dp.rf.rf_12_<7>) );
	DFFPOSX1 DFFPOSX1_105 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3166), .Q(dp.rf.rf_12_<8>) );
	DFFPOSX1 DFFPOSX1_106 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3167), .Q(dp.rf.rf_12_<9>) );
	DFFPOSX1 DFFPOSX1_107 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3168), .Q(dp.rf.rf_12_<10>) );
	DFFPOSX1 DFFPOSX1_108 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3169), .Q(dp.rf.rf_12_<11>) );
	DFFPOSX1 DFFPOSX1_109 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3170), .Q(dp.rf.rf_12_<12>) );
	DFFPOSX1 DFFPOSX1_110 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3171), .Q(dp.rf.rf_12_<13>) );
	DFFPOSX1 DFFPOSX1_111 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3172), .Q(dp.rf.rf_12_<14>) );
	DFFPOSX1 DFFPOSX1_112 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3173), .Q(dp.rf.rf_12_<15>) );
	DFFPOSX1 DFFPOSX1_113 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3174), .Q(dp.rf.rf_12_<16>) );
	DFFPOSX1 DFFPOSX1_114 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3175), .Q(dp.rf.rf_12_<17>) );
	DFFPOSX1 DFFPOSX1_115 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3176), .Q(dp.rf.rf_12_<18>) );
	DFFPOSX1 DFFPOSX1_116 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3177), .Q(dp.rf.rf_12_<19>) );
	DFFPOSX1 DFFPOSX1_117 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3178), .Q(dp.rf.rf_12_<20>) );
	DFFPOSX1 DFFPOSX1_118 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3179), .Q(dp.rf.rf_12_<21>) );
	DFFPOSX1 DFFPOSX1_119 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3180), .Q(dp.rf.rf_12_<22>) );
	DFFPOSX1 DFFPOSX1_120 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3181), .Q(dp.rf.rf_12_<23>) );
	DFFPOSX1 DFFPOSX1_121 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3182), .Q(dp.rf.rf_12_<24>) );
	DFFPOSX1 DFFPOSX1_122 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3183), .Q(dp.rf.rf_12_<25>) );
	DFFPOSX1 DFFPOSX1_123 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3184), .Q(dp.rf.rf_12_<26>) );
	DFFPOSX1 DFFPOSX1_124 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3185), .Q(dp.rf.rf_12_<27>) );
	DFFPOSX1 DFFPOSX1_125 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3186), .Q(dp.rf.rf_12_<28>) );
	DFFPOSX1 DFFPOSX1_126 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3187), .Q(dp.rf.rf_12_<29>) );
	DFFPOSX1 DFFPOSX1_127 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3188), .Q(dp.rf.rf_12_<30>) );
	DFFPOSX1 DFFPOSX1_128 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3189), .Q(dp.rf.rf_12_<31>) );
	DFFPOSX1 DFFPOSX1_129 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3190), .Q(dp.rf.rf_13_<0>) );
	DFFPOSX1 DFFPOSX1_130 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3191), .Q(dp.rf.rf_13_<1>) );
	DFFPOSX1 DFFPOSX1_131 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3192), .Q(dp.rf.rf_13_<2>) );
	DFFPOSX1 DFFPOSX1_132 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3193), .Q(dp.rf.rf_13_<3>) );
	DFFPOSX1 DFFPOSX1_133 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3194), .Q(dp.rf.rf_13_<4>) );
	DFFPOSX1 DFFPOSX1_134 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3195), .Q(dp.rf.rf_13_<5>) );
	DFFPOSX1 DFFPOSX1_135 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3196), .Q(dp.rf.rf_13_<6>) );
	DFFPOSX1 DFFPOSX1_136 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3197), .Q(dp.rf.rf_13_<7>) );
	DFFPOSX1 DFFPOSX1_137 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3198), .Q(dp.rf.rf_13_<8>) );
	DFFPOSX1 DFFPOSX1_138 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3199), .Q(dp.rf.rf_13_<9>) );
	DFFPOSX1 DFFPOSX1_139 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3200), .Q(dp.rf.rf_13_<10>) );
	DFFPOSX1 DFFPOSX1_140 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3201), .Q(dp.rf.rf_13_<11>) );
	DFFPOSX1 DFFPOSX1_141 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3202), .Q(dp.rf.rf_13_<12>) );
	DFFPOSX1 DFFPOSX1_142 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3203), .Q(dp.rf.rf_13_<13>) );
	DFFPOSX1 DFFPOSX1_143 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3204), .Q(dp.rf.rf_13_<14>) );
	DFFPOSX1 DFFPOSX1_144 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3205), .Q(dp.rf.rf_13_<15>) );
	DFFPOSX1 DFFPOSX1_145 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3206), .Q(dp.rf.rf_13_<16>) );
	DFFPOSX1 DFFPOSX1_146 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3207), .Q(dp.rf.rf_13_<17>) );
	DFFPOSX1 DFFPOSX1_147 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3208), .Q(dp.rf.rf_13_<18>) );
	DFFPOSX1 DFFPOSX1_148 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3209), .Q(dp.rf.rf_13_<19>) );
	DFFPOSX1 DFFPOSX1_149 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3210), .Q(dp.rf.rf_13_<20>) );
	DFFPOSX1 DFFPOSX1_150 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3211), .Q(dp.rf.rf_13_<21>) );
	DFFPOSX1 DFFPOSX1_151 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3212), .Q(dp.rf.rf_13_<22>) );
	DFFPOSX1 DFFPOSX1_152 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3213), .Q(dp.rf.rf_13_<23>) );
	DFFPOSX1 DFFPOSX1_153 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3214), .Q(dp.rf.rf_13_<24>) );
	DFFPOSX1 DFFPOSX1_154 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3215), .Q(dp.rf.rf_13_<25>) );
	DFFPOSX1 DFFPOSX1_155 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3216), .Q(dp.rf.rf_13_<26>) );
	DFFPOSX1 DFFPOSX1_156 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3217), .Q(dp.rf.rf_13_<27>) );
	DFFPOSX1 DFFPOSX1_157 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3218), .Q(dp.rf.rf_13_<28>) );
	DFFPOSX1 DFFPOSX1_158 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3219), .Q(dp.rf.rf_13_<29>) );
	DFFPOSX1 DFFPOSX1_159 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3220), .Q(dp.rf.rf_13_<30>) );
	DFFPOSX1 DFFPOSX1_160 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3221), .Q(dp.rf.rf_13_<31>) );
	DFFPOSX1 DFFPOSX1_161 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3222), .Q(dp.rf.rf_14_<0>) );
	DFFPOSX1 DFFPOSX1_162 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3223), .Q(dp.rf.rf_14_<1>) );
	DFFPOSX1 DFFPOSX1_163 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3224), .Q(dp.rf.rf_14_<2>) );
	DFFPOSX1 DFFPOSX1_164 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3225), .Q(dp.rf.rf_14_<3>) );
	DFFPOSX1 DFFPOSX1_165 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3226), .Q(dp.rf.rf_14_<4>) );
	DFFPOSX1 DFFPOSX1_166 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3227), .Q(dp.rf.rf_14_<5>) );
	DFFPOSX1 DFFPOSX1_167 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3228), .Q(dp.rf.rf_14_<6>) );
	DFFPOSX1 DFFPOSX1_168 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3229), .Q(dp.rf.rf_14_<7>) );
	DFFPOSX1 DFFPOSX1_169 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3230), .Q(dp.rf.rf_14_<8>) );
	DFFPOSX1 DFFPOSX1_170 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3231), .Q(dp.rf.rf_14_<9>) );
	DFFPOSX1 DFFPOSX1_171 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3232), .Q(dp.rf.rf_14_<10>) );
	DFFPOSX1 DFFPOSX1_172 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3233), .Q(dp.rf.rf_14_<11>) );
	DFFPOSX1 DFFPOSX1_173 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3234), .Q(dp.rf.rf_14_<12>) );
	DFFPOSX1 DFFPOSX1_174 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3235), .Q(dp.rf.rf_14_<13>) );
	DFFPOSX1 DFFPOSX1_175 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3236), .Q(dp.rf.rf_14_<14>) );
	DFFPOSX1 DFFPOSX1_176 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3237), .Q(dp.rf.rf_14_<15>) );
	DFFPOSX1 DFFPOSX1_177 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3238), .Q(dp.rf.rf_14_<16>) );
	DFFPOSX1 DFFPOSX1_178 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3239), .Q(dp.rf.rf_14_<17>) );
	DFFPOSX1 DFFPOSX1_179 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3240), .Q(dp.rf.rf_14_<18>) );
	DFFPOSX1 DFFPOSX1_180 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3241), .Q(dp.rf.rf_14_<19>) );
	DFFPOSX1 DFFPOSX1_181 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3242), .Q(dp.rf.rf_14_<20>) );
	DFFPOSX1 DFFPOSX1_182 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3243), .Q(dp.rf.rf_14_<21>) );
	DFFPOSX1 DFFPOSX1_183 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3244), .Q(dp.rf.rf_14_<22>) );
	DFFPOSX1 DFFPOSX1_184 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3245), .Q(dp.rf.rf_14_<23>) );
	DFFPOSX1 DFFPOSX1_185 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3246), .Q(dp.rf.rf_14_<24>) );
	DFFPOSX1 DFFPOSX1_186 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3247), .Q(dp.rf.rf_14_<25>) );
	DFFPOSX1 DFFPOSX1_187 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3248), .Q(dp.rf.rf_14_<26>) );
	DFFPOSX1 DFFPOSX1_188 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3249), .Q(dp.rf.rf_14_<27>) );
	DFFPOSX1 DFFPOSX1_189 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3250), .Q(dp.rf.rf_14_<28>) );
	DFFPOSX1 DFFPOSX1_190 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3251), .Q(dp.rf.rf_14_<29>) );
	DFFPOSX1 DFFPOSX1_191 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3252), .Q(dp.rf.rf_14_<30>) );
	DFFPOSX1 DFFPOSX1_192 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3253), .Q(dp.rf.rf_14_<31>) );
	DFFPOSX1 DFFPOSX1_193 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3254), .Q(dp.rf.rf_15_<0>) );
	DFFPOSX1 DFFPOSX1_194 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3255), .Q(dp.rf.rf_15_<1>) );
	DFFPOSX1 DFFPOSX1_195 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3256), .Q(dp.rf.rf_15_<2>) );
	DFFPOSX1 DFFPOSX1_196 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3257), .Q(dp.rf.rf_15_<3>) );
	DFFPOSX1 DFFPOSX1_197 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3258), .Q(dp.rf.rf_15_<4>) );
	DFFPOSX1 DFFPOSX1_198 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3259), .Q(dp.rf.rf_15_<5>) );
	DFFPOSX1 DFFPOSX1_199 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3260), .Q(dp.rf.rf_15_<6>) );
	DFFPOSX1 DFFPOSX1_200 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3261), .Q(dp.rf.rf_15_<7>) );
	DFFPOSX1 DFFPOSX1_201 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3262), .Q(dp.rf.rf_15_<8>) );
	DFFPOSX1 DFFPOSX1_202 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3263), .Q(dp.rf.rf_15_<9>) );
	DFFPOSX1 DFFPOSX1_203 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3264), .Q(dp.rf.rf_15_<10>) );
	DFFPOSX1 DFFPOSX1_204 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3265), .Q(dp.rf.rf_15_<11>) );
	DFFPOSX1 DFFPOSX1_205 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3266), .Q(dp.rf.rf_15_<12>) );
	DFFPOSX1 DFFPOSX1_206 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3267), .Q(dp.rf.rf_15_<13>) );
	DFFPOSX1 DFFPOSX1_207 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3268), .Q(dp.rf.rf_15_<14>) );
	DFFPOSX1 DFFPOSX1_208 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3269), .Q(dp.rf.rf_15_<15>) );
	DFFPOSX1 DFFPOSX1_209 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3270), .Q(dp.rf.rf_15_<16>) );
	DFFPOSX1 DFFPOSX1_210 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3271), .Q(dp.rf.rf_15_<17>) );
	DFFPOSX1 DFFPOSX1_211 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3272), .Q(dp.rf.rf_15_<18>) );
	DFFPOSX1 DFFPOSX1_212 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3273), .Q(dp.rf.rf_15_<19>) );
	DFFPOSX1 DFFPOSX1_213 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3274), .Q(dp.rf.rf_15_<20>) );
	DFFPOSX1 DFFPOSX1_214 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3275), .Q(dp.rf.rf_15_<21>) );
	DFFPOSX1 DFFPOSX1_215 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3276), .Q(dp.rf.rf_15_<22>) );
	DFFPOSX1 DFFPOSX1_216 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3277), .Q(dp.rf.rf_15_<23>) );
	DFFPOSX1 DFFPOSX1_217 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3278), .Q(dp.rf.rf_15_<24>) );
	DFFPOSX1 DFFPOSX1_218 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3279), .Q(dp.rf.rf_15_<25>) );
	DFFPOSX1 DFFPOSX1_219 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3280), .Q(dp.rf.rf_15_<26>) );
	DFFPOSX1 DFFPOSX1_220 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3281), .Q(dp.rf.rf_15_<27>) );
	DFFPOSX1 DFFPOSX1_221 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3282), .Q(dp.rf.rf_15_<28>) );
	DFFPOSX1 DFFPOSX1_222 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3283), .Q(dp.rf.rf_15_<29>) );
	DFFPOSX1 DFFPOSX1_223 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3284), .Q(dp.rf.rf_15_<30>) );
	DFFPOSX1 DFFPOSX1_224 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3285), .Q(dp.rf.rf_15_<31>) );
	DFFPOSX1 DFFPOSX1_225 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3286), .Q(dp.rf.rf_16_<0>) );
	DFFPOSX1 DFFPOSX1_226 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3287), .Q(dp.rf.rf_16_<1>) );
	DFFPOSX1 DFFPOSX1_227 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3288), .Q(dp.rf.rf_16_<2>) );
	DFFPOSX1 DFFPOSX1_228 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3289), .Q(dp.rf.rf_16_<3>) );
	DFFPOSX1 DFFPOSX1_229 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3290), .Q(dp.rf.rf_16_<4>) );
	DFFPOSX1 DFFPOSX1_230 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3291), .Q(dp.rf.rf_16_<5>) );
	DFFPOSX1 DFFPOSX1_231 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3292), .Q(dp.rf.rf_16_<6>) );
	DFFPOSX1 DFFPOSX1_232 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3293), .Q(dp.rf.rf_16_<7>) );
	DFFPOSX1 DFFPOSX1_233 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3294), .Q(dp.rf.rf_16_<8>) );
	DFFPOSX1 DFFPOSX1_234 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3295), .Q(dp.rf.rf_16_<9>) );
	DFFPOSX1 DFFPOSX1_235 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3296), .Q(dp.rf.rf_16_<10>) );
	DFFPOSX1 DFFPOSX1_236 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3297), .Q(dp.rf.rf_16_<11>) );
	DFFPOSX1 DFFPOSX1_237 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3298), .Q(dp.rf.rf_16_<12>) );
	DFFPOSX1 DFFPOSX1_238 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3299), .Q(dp.rf.rf_16_<13>) );
	DFFPOSX1 DFFPOSX1_239 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3300), .Q(dp.rf.rf_16_<14>) );
	DFFPOSX1 DFFPOSX1_240 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3301), .Q(dp.rf.rf_16_<15>) );
	DFFPOSX1 DFFPOSX1_241 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3302), .Q(dp.rf.rf_16_<16>) );
	DFFPOSX1 DFFPOSX1_242 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3303), .Q(dp.rf.rf_16_<17>) );
	DFFPOSX1 DFFPOSX1_243 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3304), .Q(dp.rf.rf_16_<18>) );
	DFFPOSX1 DFFPOSX1_244 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3305), .Q(dp.rf.rf_16_<19>) );
	DFFPOSX1 DFFPOSX1_245 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3306), .Q(dp.rf.rf_16_<20>) );
	DFFPOSX1 DFFPOSX1_246 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3307), .Q(dp.rf.rf_16_<21>) );
	DFFPOSX1 DFFPOSX1_247 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3308), .Q(dp.rf.rf_16_<22>) );
	DFFPOSX1 DFFPOSX1_248 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3309), .Q(dp.rf.rf_16_<23>) );
	DFFPOSX1 DFFPOSX1_249 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3310), .Q(dp.rf.rf_16_<24>) );
	DFFPOSX1 DFFPOSX1_250 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3311), .Q(dp.rf.rf_16_<25>) );
	DFFPOSX1 DFFPOSX1_251 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3312), .Q(dp.rf.rf_16_<26>) );
	DFFPOSX1 DFFPOSX1_252 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3313), .Q(dp.rf.rf_16_<27>) );
	DFFPOSX1 DFFPOSX1_253 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3314), .Q(dp.rf.rf_16_<28>) );
	DFFPOSX1 DFFPOSX1_254 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3315), .Q(dp.rf.rf_16_<29>) );
	DFFPOSX1 DFFPOSX1_255 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3316), .Q(dp.rf.rf_16_<30>) );
	DFFPOSX1 DFFPOSX1_256 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3317), .Q(dp.rf.rf_16_<31>) );
	DFFPOSX1 DFFPOSX1_257 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3318), .Q(dp.rf.rf_17_<0>) );
	DFFPOSX1 DFFPOSX1_258 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3319), .Q(dp.rf.rf_17_<1>) );
	DFFPOSX1 DFFPOSX1_259 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3320), .Q(dp.rf.rf_17_<2>) );
	DFFPOSX1 DFFPOSX1_260 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3321), .Q(dp.rf.rf_17_<3>) );
	DFFPOSX1 DFFPOSX1_261 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3322), .Q(dp.rf.rf_17_<4>) );
	DFFPOSX1 DFFPOSX1_262 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3323), .Q(dp.rf.rf_17_<5>) );
	DFFPOSX1 DFFPOSX1_263 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3324), .Q(dp.rf.rf_17_<6>) );
	DFFPOSX1 DFFPOSX1_264 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3325), .Q(dp.rf.rf_17_<7>) );
	DFFPOSX1 DFFPOSX1_265 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3326), .Q(dp.rf.rf_17_<8>) );
	DFFPOSX1 DFFPOSX1_266 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3327), .Q(dp.rf.rf_17_<9>) );
	DFFPOSX1 DFFPOSX1_267 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3328), .Q(dp.rf.rf_17_<10>) );
	DFFPOSX1 DFFPOSX1_268 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3329), .Q(dp.rf.rf_17_<11>) );
	DFFPOSX1 DFFPOSX1_269 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3330), .Q(dp.rf.rf_17_<12>) );
	DFFPOSX1 DFFPOSX1_270 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3331), .Q(dp.rf.rf_17_<13>) );
	DFFPOSX1 DFFPOSX1_271 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3332), .Q(dp.rf.rf_17_<14>) );
	DFFPOSX1 DFFPOSX1_272 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3333), .Q(dp.rf.rf_17_<15>) );
	DFFPOSX1 DFFPOSX1_273 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3334), .Q(dp.rf.rf_17_<16>) );
	DFFPOSX1 DFFPOSX1_274 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3335), .Q(dp.rf.rf_17_<17>) );
	DFFPOSX1 DFFPOSX1_275 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3336), .Q(dp.rf.rf_17_<18>) );
	DFFPOSX1 DFFPOSX1_276 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3337), .Q(dp.rf.rf_17_<19>) );
	DFFPOSX1 DFFPOSX1_277 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3338), .Q(dp.rf.rf_17_<20>) );
	DFFPOSX1 DFFPOSX1_278 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3339), .Q(dp.rf.rf_17_<21>) );
	DFFPOSX1 DFFPOSX1_279 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3340), .Q(dp.rf.rf_17_<22>) );
	DFFPOSX1 DFFPOSX1_280 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3341), .Q(dp.rf.rf_17_<23>) );
	DFFPOSX1 DFFPOSX1_281 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3342), .Q(dp.rf.rf_17_<24>) );
	DFFPOSX1 DFFPOSX1_282 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3343), .Q(dp.rf.rf_17_<25>) );
	DFFPOSX1 DFFPOSX1_283 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3344), .Q(dp.rf.rf_17_<26>) );
	DFFPOSX1 DFFPOSX1_284 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3345), .Q(dp.rf.rf_17_<27>) );
	DFFPOSX1 DFFPOSX1_285 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3346), .Q(dp.rf.rf_17_<28>) );
	DFFPOSX1 DFFPOSX1_286 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3347), .Q(dp.rf.rf_17_<29>) );
	DFFPOSX1 DFFPOSX1_287 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3348), .Q(dp.rf.rf_17_<30>) );
	DFFPOSX1 DFFPOSX1_288 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3349), .Q(dp.rf.rf_17_<31>) );
	DFFPOSX1 DFFPOSX1_289 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3350), .Q(dp.rf.rf_18_<0>) );
	DFFPOSX1 DFFPOSX1_290 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3351), .Q(dp.rf.rf_18_<1>) );
	DFFPOSX1 DFFPOSX1_291 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3352), .Q(dp.rf.rf_18_<2>) );
	DFFPOSX1 DFFPOSX1_292 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3353), .Q(dp.rf.rf_18_<3>) );
	DFFPOSX1 DFFPOSX1_293 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3354), .Q(dp.rf.rf_18_<4>) );
	DFFPOSX1 DFFPOSX1_294 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3355), .Q(dp.rf.rf_18_<5>) );
	DFFPOSX1 DFFPOSX1_295 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3356), .Q(dp.rf.rf_18_<6>) );
	DFFPOSX1 DFFPOSX1_296 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3357), .Q(dp.rf.rf_18_<7>) );
	DFFPOSX1 DFFPOSX1_297 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3358), .Q(dp.rf.rf_18_<8>) );
	DFFPOSX1 DFFPOSX1_298 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3359), .Q(dp.rf.rf_18_<9>) );
	DFFPOSX1 DFFPOSX1_299 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3360), .Q(dp.rf.rf_18_<10>) );
	DFFPOSX1 DFFPOSX1_300 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3361), .Q(dp.rf.rf_18_<11>) );
	DFFPOSX1 DFFPOSX1_301 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3362), .Q(dp.rf.rf_18_<12>) );
	DFFPOSX1 DFFPOSX1_302 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3363), .Q(dp.rf.rf_18_<13>) );
	DFFPOSX1 DFFPOSX1_303 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3364), .Q(dp.rf.rf_18_<14>) );
	DFFPOSX1 DFFPOSX1_304 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3365), .Q(dp.rf.rf_18_<15>) );
	DFFPOSX1 DFFPOSX1_305 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3366), .Q(dp.rf.rf_18_<16>) );
	DFFPOSX1 DFFPOSX1_306 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3367), .Q(dp.rf.rf_18_<17>) );
	DFFPOSX1 DFFPOSX1_307 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3368), .Q(dp.rf.rf_18_<18>) );
	DFFPOSX1 DFFPOSX1_308 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3369), .Q(dp.rf.rf_18_<19>) );
	DFFPOSX1 DFFPOSX1_309 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3370), .Q(dp.rf.rf_18_<20>) );
	DFFPOSX1 DFFPOSX1_310 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3371), .Q(dp.rf.rf_18_<21>) );
	DFFPOSX1 DFFPOSX1_311 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3372), .Q(dp.rf.rf_18_<22>) );
	DFFPOSX1 DFFPOSX1_312 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3373), .Q(dp.rf.rf_18_<23>) );
	DFFPOSX1 DFFPOSX1_313 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3374), .Q(dp.rf.rf_18_<24>) );
	DFFPOSX1 DFFPOSX1_314 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3375), .Q(dp.rf.rf_18_<25>) );
	DFFPOSX1 DFFPOSX1_315 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3376), .Q(dp.rf.rf_18_<26>) );
	DFFPOSX1 DFFPOSX1_316 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3377), .Q(dp.rf.rf_18_<27>) );
	DFFPOSX1 DFFPOSX1_317 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3378), .Q(dp.rf.rf_18_<28>) );
	DFFPOSX1 DFFPOSX1_318 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3379), .Q(dp.rf.rf_18_<29>) );
	DFFPOSX1 DFFPOSX1_319 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3380), .Q(dp.rf.rf_18_<30>) );
	DFFPOSX1 DFFPOSX1_320 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3381), .Q(dp.rf.rf_18_<31>) );
	DFFPOSX1 DFFPOSX1_321 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3382), .Q(dp.rf.rf_19_<0>) );
	DFFPOSX1 DFFPOSX1_322 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3383), .Q(dp.rf.rf_19_<1>) );
	DFFPOSX1 DFFPOSX1_323 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3384), .Q(dp.rf.rf_19_<2>) );
	DFFPOSX1 DFFPOSX1_324 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3385), .Q(dp.rf.rf_19_<3>) );
	DFFPOSX1 DFFPOSX1_325 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3386), .Q(dp.rf.rf_19_<4>) );
	DFFPOSX1 DFFPOSX1_326 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3387), .Q(dp.rf.rf_19_<5>) );
	DFFPOSX1 DFFPOSX1_327 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3388), .Q(dp.rf.rf_19_<6>) );
	DFFPOSX1 DFFPOSX1_328 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3389), .Q(dp.rf.rf_19_<7>) );
	DFFPOSX1 DFFPOSX1_329 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3390), .Q(dp.rf.rf_19_<8>) );
	DFFPOSX1 DFFPOSX1_330 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3391), .Q(dp.rf.rf_19_<9>) );
	DFFPOSX1 DFFPOSX1_331 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3392), .Q(dp.rf.rf_19_<10>) );
	DFFPOSX1 DFFPOSX1_332 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3393), .Q(dp.rf.rf_19_<11>) );
	DFFPOSX1 DFFPOSX1_333 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3394), .Q(dp.rf.rf_19_<12>) );
	DFFPOSX1 DFFPOSX1_334 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3395), .Q(dp.rf.rf_19_<13>) );
	DFFPOSX1 DFFPOSX1_335 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3396), .Q(dp.rf.rf_19_<14>) );
	DFFPOSX1 DFFPOSX1_336 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3397), .Q(dp.rf.rf_19_<15>) );
	DFFPOSX1 DFFPOSX1_337 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3398), .Q(dp.rf.rf_19_<16>) );
	DFFPOSX1 DFFPOSX1_338 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3399), .Q(dp.rf.rf_19_<17>) );
	DFFPOSX1 DFFPOSX1_339 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3400), .Q(dp.rf.rf_19_<18>) );
	DFFPOSX1 DFFPOSX1_340 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3401), .Q(dp.rf.rf_19_<19>) );
	DFFPOSX1 DFFPOSX1_341 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3402), .Q(dp.rf.rf_19_<20>) );
	DFFPOSX1 DFFPOSX1_342 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3403), .Q(dp.rf.rf_19_<21>) );
	DFFPOSX1 DFFPOSX1_343 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3404), .Q(dp.rf.rf_19_<22>) );
	DFFPOSX1 DFFPOSX1_344 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3405), .Q(dp.rf.rf_19_<23>) );
	DFFPOSX1 DFFPOSX1_345 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3406), .Q(dp.rf.rf_19_<24>) );
	DFFPOSX1 DFFPOSX1_346 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3407), .Q(dp.rf.rf_19_<25>) );
	DFFPOSX1 DFFPOSX1_347 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3408), .Q(dp.rf.rf_19_<26>) );
	DFFPOSX1 DFFPOSX1_348 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3409), .Q(dp.rf.rf_19_<27>) );
	DFFPOSX1 DFFPOSX1_349 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3410), .Q(dp.rf.rf_19_<28>) );
	DFFPOSX1 DFFPOSX1_350 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3411), .Q(dp.rf.rf_19_<29>) );
	DFFPOSX1 DFFPOSX1_351 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3412), .Q(dp.rf.rf_19_<30>) );
	DFFPOSX1 DFFPOSX1_352 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3413), .Q(dp.rf.rf_19_<31>) );
	DFFPOSX1 DFFPOSX1_353 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3414), .Q(dp.rf.rf_1_<0>) );
	DFFPOSX1 DFFPOSX1_354 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3415), .Q(dp.rf.rf_1_<1>) );
	DFFPOSX1 DFFPOSX1_355 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3416), .Q(dp.rf.rf_1_<2>) );
	DFFPOSX1 DFFPOSX1_356 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3417), .Q(dp.rf.rf_1_<3>) );
	DFFPOSX1 DFFPOSX1_357 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3418), .Q(dp.rf.rf_1_<4>) );
	DFFPOSX1 DFFPOSX1_358 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3419), .Q(dp.rf.rf_1_<5>) );
	DFFPOSX1 DFFPOSX1_359 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3420), .Q(dp.rf.rf_1_<6>) );
	DFFPOSX1 DFFPOSX1_360 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3421), .Q(dp.rf.rf_1_<7>) );
	DFFPOSX1 DFFPOSX1_361 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3422), .Q(dp.rf.rf_1_<8>) );
	DFFPOSX1 DFFPOSX1_362 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3423), .Q(dp.rf.rf_1_<9>) );
	DFFPOSX1 DFFPOSX1_363 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3424), .Q(dp.rf.rf_1_<10>) );
	DFFPOSX1 DFFPOSX1_364 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3425), .Q(dp.rf.rf_1_<11>) );
	DFFPOSX1 DFFPOSX1_365 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3426), .Q(dp.rf.rf_1_<12>) );
	DFFPOSX1 DFFPOSX1_366 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3427), .Q(dp.rf.rf_1_<13>) );
	DFFPOSX1 DFFPOSX1_367 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3428), .Q(dp.rf.rf_1_<14>) );
	DFFPOSX1 DFFPOSX1_368 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3429), .Q(dp.rf.rf_1_<15>) );
	DFFPOSX1 DFFPOSX1_369 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3430), .Q(dp.rf.rf_1_<16>) );
	DFFPOSX1 DFFPOSX1_370 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3431), .Q(dp.rf.rf_1_<17>) );
	DFFPOSX1 DFFPOSX1_371 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3432), .Q(dp.rf.rf_1_<18>) );
	DFFPOSX1 DFFPOSX1_372 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3433), .Q(dp.rf.rf_1_<19>) );
	DFFPOSX1 DFFPOSX1_373 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3434), .Q(dp.rf.rf_1_<20>) );
	DFFPOSX1 DFFPOSX1_374 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3435), .Q(dp.rf.rf_1_<21>) );
	DFFPOSX1 DFFPOSX1_375 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3436), .Q(dp.rf.rf_1_<22>) );
	DFFPOSX1 DFFPOSX1_376 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3437), .Q(dp.rf.rf_1_<23>) );
	DFFPOSX1 DFFPOSX1_377 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3438), .Q(dp.rf.rf_1_<24>) );
	DFFPOSX1 DFFPOSX1_378 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3439), .Q(dp.rf.rf_1_<25>) );
	DFFPOSX1 DFFPOSX1_379 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3440), .Q(dp.rf.rf_1_<26>) );
	DFFPOSX1 DFFPOSX1_380 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3441), .Q(dp.rf.rf_1_<27>) );
	DFFPOSX1 DFFPOSX1_381 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3442), .Q(dp.rf.rf_1_<28>) );
	DFFPOSX1 DFFPOSX1_382 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3443), .Q(dp.rf.rf_1_<29>) );
	DFFPOSX1 DFFPOSX1_383 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3444), .Q(dp.rf.rf_1_<30>) );
	DFFPOSX1 DFFPOSX1_384 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3445), .Q(dp.rf.rf_1_<31>) );
	DFFPOSX1 DFFPOSX1_385 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3446), .Q(dp.rf.rf_20_<0>) );
	DFFPOSX1 DFFPOSX1_386 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3447), .Q(dp.rf.rf_20_<1>) );
	DFFPOSX1 DFFPOSX1_387 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3448), .Q(dp.rf.rf_20_<2>) );
	DFFPOSX1 DFFPOSX1_388 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3449), .Q(dp.rf.rf_20_<3>) );
	DFFPOSX1 DFFPOSX1_389 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3450), .Q(dp.rf.rf_20_<4>) );
	DFFPOSX1 DFFPOSX1_390 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3451), .Q(dp.rf.rf_20_<5>) );
	DFFPOSX1 DFFPOSX1_391 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3452), .Q(dp.rf.rf_20_<6>) );
	DFFPOSX1 DFFPOSX1_392 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3453), .Q(dp.rf.rf_20_<7>) );
	DFFPOSX1 DFFPOSX1_393 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3454), .Q(dp.rf.rf_20_<8>) );
	DFFPOSX1 DFFPOSX1_394 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3455), .Q(dp.rf.rf_20_<9>) );
	DFFPOSX1 DFFPOSX1_395 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3456), .Q(dp.rf.rf_20_<10>) );
	DFFPOSX1 DFFPOSX1_396 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3457), .Q(dp.rf.rf_20_<11>) );
	DFFPOSX1 DFFPOSX1_397 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3458), .Q(dp.rf.rf_20_<12>) );
	DFFPOSX1 DFFPOSX1_398 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3459), .Q(dp.rf.rf_20_<13>) );
	DFFPOSX1 DFFPOSX1_399 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3460), .Q(dp.rf.rf_20_<14>) );
	DFFPOSX1 DFFPOSX1_400 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3461), .Q(dp.rf.rf_20_<15>) );
	DFFPOSX1 DFFPOSX1_401 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3462), .Q(dp.rf.rf_20_<16>) );
	DFFPOSX1 DFFPOSX1_402 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3463), .Q(dp.rf.rf_20_<17>) );
	DFFPOSX1 DFFPOSX1_403 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3464), .Q(dp.rf.rf_20_<18>) );
	DFFPOSX1 DFFPOSX1_404 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3465), .Q(dp.rf.rf_20_<19>) );
	DFFPOSX1 DFFPOSX1_405 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3466), .Q(dp.rf.rf_20_<20>) );
	DFFPOSX1 DFFPOSX1_406 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3467), .Q(dp.rf.rf_20_<21>) );
	DFFPOSX1 DFFPOSX1_407 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3468), .Q(dp.rf.rf_20_<22>) );
	DFFPOSX1 DFFPOSX1_408 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3469), .Q(dp.rf.rf_20_<23>) );
	DFFPOSX1 DFFPOSX1_409 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3470), .Q(dp.rf.rf_20_<24>) );
	DFFPOSX1 DFFPOSX1_410 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3471), .Q(dp.rf.rf_20_<25>) );
	DFFPOSX1 DFFPOSX1_411 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3472), .Q(dp.rf.rf_20_<26>) );
	DFFPOSX1 DFFPOSX1_412 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3473), .Q(dp.rf.rf_20_<27>) );
	DFFPOSX1 DFFPOSX1_413 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3474), .Q(dp.rf.rf_20_<28>) );
	DFFPOSX1 DFFPOSX1_414 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3475), .Q(dp.rf.rf_20_<29>) );
	DFFPOSX1 DFFPOSX1_415 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3476), .Q(dp.rf.rf_20_<30>) );
	DFFPOSX1 DFFPOSX1_416 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3477), .Q(dp.rf.rf_20_<31>) );
	DFFPOSX1 DFFPOSX1_417 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3478), .Q(dp.rf.rf_21_<0>) );
	DFFPOSX1 DFFPOSX1_418 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3479), .Q(dp.rf.rf_21_<1>) );
	DFFPOSX1 DFFPOSX1_419 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3480), .Q(dp.rf.rf_21_<2>) );
	DFFPOSX1 DFFPOSX1_420 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3481), .Q(dp.rf.rf_21_<3>) );
	DFFPOSX1 DFFPOSX1_421 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3482), .Q(dp.rf.rf_21_<4>) );
	DFFPOSX1 DFFPOSX1_422 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3483), .Q(dp.rf.rf_21_<5>) );
	DFFPOSX1 DFFPOSX1_423 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3484), .Q(dp.rf.rf_21_<6>) );
	DFFPOSX1 DFFPOSX1_424 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3485), .Q(dp.rf.rf_21_<7>) );
	DFFPOSX1 DFFPOSX1_425 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3486), .Q(dp.rf.rf_21_<8>) );
	DFFPOSX1 DFFPOSX1_426 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3487), .Q(dp.rf.rf_21_<9>) );
	DFFPOSX1 DFFPOSX1_427 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3488), .Q(dp.rf.rf_21_<10>) );
	DFFPOSX1 DFFPOSX1_428 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3489), .Q(dp.rf.rf_21_<11>) );
	DFFPOSX1 DFFPOSX1_429 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3490), .Q(dp.rf.rf_21_<12>) );
	DFFPOSX1 DFFPOSX1_430 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3491), .Q(dp.rf.rf_21_<13>) );
	DFFPOSX1 DFFPOSX1_431 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3492), .Q(dp.rf.rf_21_<14>) );
	DFFPOSX1 DFFPOSX1_432 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3493), .Q(dp.rf.rf_21_<15>) );
	DFFPOSX1 DFFPOSX1_433 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3494), .Q(dp.rf.rf_21_<16>) );
	DFFPOSX1 DFFPOSX1_434 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3495), .Q(dp.rf.rf_21_<17>) );
	DFFPOSX1 DFFPOSX1_435 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3496), .Q(dp.rf.rf_21_<18>) );
	DFFPOSX1 DFFPOSX1_436 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3497), .Q(dp.rf.rf_21_<19>) );
	DFFPOSX1 DFFPOSX1_437 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3498), .Q(dp.rf.rf_21_<20>) );
	DFFPOSX1 DFFPOSX1_438 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3499), .Q(dp.rf.rf_21_<21>) );
	DFFPOSX1 DFFPOSX1_439 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3500), .Q(dp.rf.rf_21_<22>) );
	DFFPOSX1 DFFPOSX1_440 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3501), .Q(dp.rf.rf_21_<23>) );
	DFFPOSX1 DFFPOSX1_441 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3502), .Q(dp.rf.rf_21_<24>) );
	DFFPOSX1 DFFPOSX1_442 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3503), .Q(dp.rf.rf_21_<25>) );
	DFFPOSX1 DFFPOSX1_443 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3504), .Q(dp.rf.rf_21_<26>) );
	DFFPOSX1 DFFPOSX1_444 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3505), .Q(dp.rf.rf_21_<27>) );
	DFFPOSX1 DFFPOSX1_445 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3506), .Q(dp.rf.rf_21_<28>) );
	DFFPOSX1 DFFPOSX1_446 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3507), .Q(dp.rf.rf_21_<29>) );
	DFFPOSX1 DFFPOSX1_447 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3508), .Q(dp.rf.rf_21_<30>) );
	DFFPOSX1 DFFPOSX1_448 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3509), .Q(dp.rf.rf_21_<31>) );
	DFFPOSX1 DFFPOSX1_449 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3510), .Q(dp.rf.rf_22_<0>) );
	DFFPOSX1 DFFPOSX1_450 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3511), .Q(dp.rf.rf_22_<1>) );
	DFFPOSX1 DFFPOSX1_451 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3512), .Q(dp.rf.rf_22_<2>) );
	DFFPOSX1 DFFPOSX1_452 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3513), .Q(dp.rf.rf_22_<3>) );
	DFFPOSX1 DFFPOSX1_453 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3514), .Q(dp.rf.rf_22_<4>) );
	DFFPOSX1 DFFPOSX1_454 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3515), .Q(dp.rf.rf_22_<5>) );
	DFFPOSX1 DFFPOSX1_455 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3516), .Q(dp.rf.rf_22_<6>) );
	DFFPOSX1 DFFPOSX1_456 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3517), .Q(dp.rf.rf_22_<7>) );
	DFFPOSX1 DFFPOSX1_457 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3518), .Q(dp.rf.rf_22_<8>) );
	DFFPOSX1 DFFPOSX1_458 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3519), .Q(dp.rf.rf_22_<9>) );
	DFFPOSX1 DFFPOSX1_459 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3520), .Q(dp.rf.rf_22_<10>) );
	DFFPOSX1 DFFPOSX1_460 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3521), .Q(dp.rf.rf_22_<11>) );
	DFFPOSX1 DFFPOSX1_461 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3522), .Q(dp.rf.rf_22_<12>) );
	DFFPOSX1 DFFPOSX1_462 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3523), .Q(dp.rf.rf_22_<13>) );
	DFFPOSX1 DFFPOSX1_463 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3524), .Q(dp.rf.rf_22_<14>) );
	DFFPOSX1 DFFPOSX1_464 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3525), .Q(dp.rf.rf_22_<15>) );
	DFFPOSX1 DFFPOSX1_465 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3526), .Q(dp.rf.rf_22_<16>) );
	DFFPOSX1 DFFPOSX1_466 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3527), .Q(dp.rf.rf_22_<17>) );
	DFFPOSX1 DFFPOSX1_467 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3528), .Q(dp.rf.rf_22_<18>) );
	DFFPOSX1 DFFPOSX1_468 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3529), .Q(dp.rf.rf_22_<19>) );
	DFFPOSX1 DFFPOSX1_469 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3530), .Q(dp.rf.rf_22_<20>) );
	DFFPOSX1 DFFPOSX1_470 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3531), .Q(dp.rf.rf_22_<21>) );
	DFFPOSX1 DFFPOSX1_471 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3532), .Q(dp.rf.rf_22_<22>) );
	DFFPOSX1 DFFPOSX1_472 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3533), .Q(dp.rf.rf_22_<23>) );
	DFFPOSX1 DFFPOSX1_473 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3534), .Q(dp.rf.rf_22_<24>) );
	DFFPOSX1 DFFPOSX1_474 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3535), .Q(dp.rf.rf_22_<25>) );
	DFFPOSX1 DFFPOSX1_475 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3536), .Q(dp.rf.rf_22_<26>) );
	DFFPOSX1 DFFPOSX1_476 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3537), .Q(dp.rf.rf_22_<27>) );
	DFFPOSX1 DFFPOSX1_477 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3538), .Q(dp.rf.rf_22_<28>) );
	DFFPOSX1 DFFPOSX1_478 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3539), .Q(dp.rf.rf_22_<29>) );
	DFFPOSX1 DFFPOSX1_479 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3540), .Q(dp.rf.rf_22_<30>) );
	DFFPOSX1 DFFPOSX1_480 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3541), .Q(dp.rf.rf_22_<31>) );
	DFFPOSX1 DFFPOSX1_481 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3542), .Q(dp.rf.rf_23_<0>) );
	DFFPOSX1 DFFPOSX1_482 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3543), .Q(dp.rf.rf_23_<1>) );
	DFFPOSX1 DFFPOSX1_483 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3544), .Q(dp.rf.rf_23_<2>) );
	DFFPOSX1 DFFPOSX1_484 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3545), .Q(dp.rf.rf_23_<3>) );
	DFFPOSX1 DFFPOSX1_485 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3546), .Q(dp.rf.rf_23_<4>) );
	DFFPOSX1 DFFPOSX1_486 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3547), .Q(dp.rf.rf_23_<5>) );
	DFFPOSX1 DFFPOSX1_487 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3548), .Q(dp.rf.rf_23_<6>) );
	DFFPOSX1 DFFPOSX1_488 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3549), .Q(dp.rf.rf_23_<7>) );
	DFFPOSX1 DFFPOSX1_489 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3550), .Q(dp.rf.rf_23_<8>) );
	DFFPOSX1 DFFPOSX1_490 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3551), .Q(dp.rf.rf_23_<9>) );
	DFFPOSX1 DFFPOSX1_491 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3552), .Q(dp.rf.rf_23_<10>) );
	DFFPOSX1 DFFPOSX1_492 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3553), .Q(dp.rf.rf_23_<11>) );
	DFFPOSX1 DFFPOSX1_493 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3554), .Q(dp.rf.rf_23_<12>) );
	DFFPOSX1 DFFPOSX1_494 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3555), .Q(dp.rf.rf_23_<13>) );
	DFFPOSX1 DFFPOSX1_495 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3556), .Q(dp.rf.rf_23_<14>) );
	DFFPOSX1 DFFPOSX1_496 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3557), .Q(dp.rf.rf_23_<15>) );
	DFFPOSX1 DFFPOSX1_497 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3558), .Q(dp.rf.rf_23_<16>) );
	DFFPOSX1 DFFPOSX1_498 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3559), .Q(dp.rf.rf_23_<17>) );
	DFFPOSX1 DFFPOSX1_499 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3560), .Q(dp.rf.rf_23_<18>) );
	DFFPOSX1 DFFPOSX1_500 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3561), .Q(dp.rf.rf_23_<19>) );
	DFFPOSX1 DFFPOSX1_501 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3562), .Q(dp.rf.rf_23_<20>) );
	DFFPOSX1 DFFPOSX1_502 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3563), .Q(dp.rf.rf_23_<21>) );
	DFFPOSX1 DFFPOSX1_503 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3564), .Q(dp.rf.rf_23_<22>) );
	DFFPOSX1 DFFPOSX1_504 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3565), .Q(dp.rf.rf_23_<23>) );
	DFFPOSX1 DFFPOSX1_505 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3566), .Q(dp.rf.rf_23_<24>) );
	DFFPOSX1 DFFPOSX1_506 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3567), .Q(dp.rf.rf_23_<25>) );
	DFFPOSX1 DFFPOSX1_507 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3568), .Q(dp.rf.rf_23_<26>) );
	DFFPOSX1 DFFPOSX1_508 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3569), .Q(dp.rf.rf_23_<27>) );
	DFFPOSX1 DFFPOSX1_509 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3570), .Q(dp.rf.rf_23_<28>) );
	DFFPOSX1 DFFPOSX1_510 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3571), .Q(dp.rf.rf_23_<29>) );
	DFFPOSX1 DFFPOSX1_511 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3572), .Q(dp.rf.rf_23_<30>) );
	DFFPOSX1 DFFPOSX1_512 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3573), .Q(dp.rf.rf_23_<31>) );
	DFFPOSX1 DFFPOSX1_513 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3574), .Q(dp.rf.rf_24_<0>) );
	DFFPOSX1 DFFPOSX1_514 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3575), .Q(dp.rf.rf_24_<1>) );
	DFFPOSX1 DFFPOSX1_515 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3576), .Q(dp.rf.rf_24_<2>) );
	DFFPOSX1 DFFPOSX1_516 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3577), .Q(dp.rf.rf_24_<3>) );
	DFFPOSX1 DFFPOSX1_517 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3578), .Q(dp.rf.rf_24_<4>) );
	DFFPOSX1 DFFPOSX1_518 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3579), .Q(dp.rf.rf_24_<5>) );
	DFFPOSX1 DFFPOSX1_519 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3580), .Q(dp.rf.rf_24_<6>) );
	DFFPOSX1 DFFPOSX1_520 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3581), .Q(dp.rf.rf_24_<7>) );
	DFFPOSX1 DFFPOSX1_521 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3582), .Q(dp.rf.rf_24_<8>) );
	DFFPOSX1 DFFPOSX1_522 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3583), .Q(dp.rf.rf_24_<9>) );
	DFFPOSX1 DFFPOSX1_523 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3584), .Q(dp.rf.rf_24_<10>) );
	DFFPOSX1 DFFPOSX1_524 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3585), .Q(dp.rf.rf_24_<11>) );
	DFFPOSX1 DFFPOSX1_525 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3586), .Q(dp.rf.rf_24_<12>) );
	DFFPOSX1 DFFPOSX1_526 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3587), .Q(dp.rf.rf_24_<13>) );
	DFFPOSX1 DFFPOSX1_527 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3588), .Q(dp.rf.rf_24_<14>) );
	DFFPOSX1 DFFPOSX1_528 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3589), .Q(dp.rf.rf_24_<15>) );
	DFFPOSX1 DFFPOSX1_529 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3590), .Q(dp.rf.rf_24_<16>) );
	DFFPOSX1 DFFPOSX1_530 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3591), .Q(dp.rf.rf_24_<17>) );
	DFFPOSX1 DFFPOSX1_531 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3592), .Q(dp.rf.rf_24_<18>) );
	DFFPOSX1 DFFPOSX1_532 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3593), .Q(dp.rf.rf_24_<19>) );
	DFFPOSX1 DFFPOSX1_533 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3594), .Q(dp.rf.rf_24_<20>) );
	DFFPOSX1 DFFPOSX1_534 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3595), .Q(dp.rf.rf_24_<21>) );
	DFFPOSX1 DFFPOSX1_535 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3596), .Q(dp.rf.rf_24_<22>) );
	DFFPOSX1 DFFPOSX1_536 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3597), .Q(dp.rf.rf_24_<23>) );
	DFFPOSX1 DFFPOSX1_537 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3598), .Q(dp.rf.rf_24_<24>) );
	DFFPOSX1 DFFPOSX1_538 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3599), .Q(dp.rf.rf_24_<25>) );
	DFFPOSX1 DFFPOSX1_539 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3600), .Q(dp.rf.rf_24_<26>) );
	DFFPOSX1 DFFPOSX1_540 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3601), .Q(dp.rf.rf_24_<27>) );
	DFFPOSX1 DFFPOSX1_541 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3602), .Q(dp.rf.rf_24_<28>) );
	DFFPOSX1 DFFPOSX1_542 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3603), .Q(dp.rf.rf_24_<29>) );
	DFFPOSX1 DFFPOSX1_543 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3604), .Q(dp.rf.rf_24_<30>) );
	DFFPOSX1 DFFPOSX1_544 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3605), .Q(dp.rf.rf_24_<31>) );
	DFFPOSX1 DFFPOSX1_545 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3606), .Q(dp.rf.rf_25_<0>) );
	DFFPOSX1 DFFPOSX1_546 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3607), .Q(dp.rf.rf_25_<1>) );
	DFFPOSX1 DFFPOSX1_547 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3608), .Q(dp.rf.rf_25_<2>) );
	DFFPOSX1 DFFPOSX1_548 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3609), .Q(dp.rf.rf_25_<3>) );
	DFFPOSX1 DFFPOSX1_549 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3610), .Q(dp.rf.rf_25_<4>) );
	DFFPOSX1 DFFPOSX1_550 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3611), .Q(dp.rf.rf_25_<5>) );
	DFFPOSX1 DFFPOSX1_551 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3612), .Q(dp.rf.rf_25_<6>) );
	DFFPOSX1 DFFPOSX1_552 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3613), .Q(dp.rf.rf_25_<7>) );
	DFFPOSX1 DFFPOSX1_553 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3614), .Q(dp.rf.rf_25_<8>) );
	DFFPOSX1 DFFPOSX1_554 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3615), .Q(dp.rf.rf_25_<9>) );
	DFFPOSX1 DFFPOSX1_555 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3616), .Q(dp.rf.rf_25_<10>) );
	DFFPOSX1 DFFPOSX1_556 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3617), .Q(dp.rf.rf_25_<11>) );
	DFFPOSX1 DFFPOSX1_557 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3618), .Q(dp.rf.rf_25_<12>) );
	DFFPOSX1 DFFPOSX1_558 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3619), .Q(dp.rf.rf_25_<13>) );
	DFFPOSX1 DFFPOSX1_559 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3620), .Q(dp.rf.rf_25_<14>) );
	DFFPOSX1 DFFPOSX1_560 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3621), .Q(dp.rf.rf_25_<15>) );
	DFFPOSX1 DFFPOSX1_561 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3622), .Q(dp.rf.rf_25_<16>) );
	DFFPOSX1 DFFPOSX1_562 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3623), .Q(dp.rf.rf_25_<17>) );
	DFFPOSX1 DFFPOSX1_563 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3624), .Q(dp.rf.rf_25_<18>) );
	DFFPOSX1 DFFPOSX1_564 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3625), .Q(dp.rf.rf_25_<19>) );
	DFFPOSX1 DFFPOSX1_565 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3626), .Q(dp.rf.rf_25_<20>) );
	DFFPOSX1 DFFPOSX1_566 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3627), .Q(dp.rf.rf_25_<21>) );
	DFFPOSX1 DFFPOSX1_567 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3628), .Q(dp.rf.rf_25_<22>) );
	DFFPOSX1 DFFPOSX1_568 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3629), .Q(dp.rf.rf_25_<23>) );
	DFFPOSX1 DFFPOSX1_569 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3630), .Q(dp.rf.rf_25_<24>) );
	DFFPOSX1 DFFPOSX1_570 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3631), .Q(dp.rf.rf_25_<25>) );
	DFFPOSX1 DFFPOSX1_571 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3632), .Q(dp.rf.rf_25_<26>) );
	DFFPOSX1 DFFPOSX1_572 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3633), .Q(dp.rf.rf_25_<27>) );
	DFFPOSX1 DFFPOSX1_573 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3634), .Q(dp.rf.rf_25_<28>) );
	DFFPOSX1 DFFPOSX1_574 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3635), .Q(dp.rf.rf_25_<29>) );
	DFFPOSX1 DFFPOSX1_575 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3636), .Q(dp.rf.rf_25_<30>) );
	DFFPOSX1 DFFPOSX1_576 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3637), .Q(dp.rf.rf_25_<31>) );
	DFFPOSX1 DFFPOSX1_577 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3638), .Q(dp.rf.rf_26_<0>) );
	DFFPOSX1 DFFPOSX1_578 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3639), .Q(dp.rf.rf_26_<1>) );
	DFFPOSX1 DFFPOSX1_579 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3640), .Q(dp.rf.rf_26_<2>) );
	DFFPOSX1 DFFPOSX1_580 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3641), .Q(dp.rf.rf_26_<3>) );
	DFFPOSX1 DFFPOSX1_581 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3642), .Q(dp.rf.rf_26_<4>) );
	DFFPOSX1 DFFPOSX1_582 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3643), .Q(dp.rf.rf_26_<5>) );
	DFFPOSX1 DFFPOSX1_583 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3644), .Q(dp.rf.rf_26_<6>) );
	DFFPOSX1 DFFPOSX1_584 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3645), .Q(dp.rf.rf_26_<7>) );
	DFFPOSX1 DFFPOSX1_585 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3646), .Q(dp.rf.rf_26_<8>) );
	DFFPOSX1 DFFPOSX1_586 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3647), .Q(dp.rf.rf_26_<9>) );
	DFFPOSX1 DFFPOSX1_587 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3648), .Q(dp.rf.rf_26_<10>) );
	DFFPOSX1 DFFPOSX1_588 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3649), .Q(dp.rf.rf_26_<11>) );
	DFFPOSX1 DFFPOSX1_589 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3650), .Q(dp.rf.rf_26_<12>) );
	DFFPOSX1 DFFPOSX1_590 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3651), .Q(dp.rf.rf_26_<13>) );
	DFFPOSX1 DFFPOSX1_591 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3652), .Q(dp.rf.rf_26_<14>) );
	DFFPOSX1 DFFPOSX1_592 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3653), .Q(dp.rf.rf_26_<15>) );
	DFFPOSX1 DFFPOSX1_593 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3654), .Q(dp.rf.rf_26_<16>) );
	DFFPOSX1 DFFPOSX1_594 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3655), .Q(dp.rf.rf_26_<17>) );
	DFFPOSX1 DFFPOSX1_595 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3656), .Q(dp.rf.rf_26_<18>) );
	DFFPOSX1 DFFPOSX1_596 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3657), .Q(dp.rf.rf_26_<19>) );
	DFFPOSX1 DFFPOSX1_597 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3658), .Q(dp.rf.rf_26_<20>) );
	DFFPOSX1 DFFPOSX1_598 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3659), .Q(dp.rf.rf_26_<21>) );
	DFFPOSX1 DFFPOSX1_599 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3660), .Q(dp.rf.rf_26_<22>) );
	DFFPOSX1 DFFPOSX1_600 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3661), .Q(dp.rf.rf_26_<23>) );
	DFFPOSX1 DFFPOSX1_601 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3662), .Q(dp.rf.rf_26_<24>) );
	DFFPOSX1 DFFPOSX1_602 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3663), .Q(dp.rf.rf_26_<25>) );
	DFFPOSX1 DFFPOSX1_603 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3664), .Q(dp.rf.rf_26_<26>) );
	DFFPOSX1 DFFPOSX1_604 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3665), .Q(dp.rf.rf_26_<27>) );
	DFFPOSX1 DFFPOSX1_605 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3666), .Q(dp.rf.rf_26_<28>) );
	DFFPOSX1 DFFPOSX1_606 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3667), .Q(dp.rf.rf_26_<29>) );
	DFFPOSX1 DFFPOSX1_607 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3668), .Q(dp.rf.rf_26_<30>) );
	DFFPOSX1 DFFPOSX1_608 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3669), .Q(dp.rf.rf_26_<31>) );
	DFFPOSX1 DFFPOSX1_609 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3670), .Q(dp.rf.rf_27_<0>) );
	DFFPOSX1 DFFPOSX1_610 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3671), .Q(dp.rf.rf_27_<1>) );
	DFFPOSX1 DFFPOSX1_611 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3672), .Q(dp.rf.rf_27_<2>) );
	DFFPOSX1 DFFPOSX1_612 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3673), .Q(dp.rf.rf_27_<3>) );
	DFFPOSX1 DFFPOSX1_613 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3674), .Q(dp.rf.rf_27_<4>) );
	DFFPOSX1 DFFPOSX1_614 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3675), .Q(dp.rf.rf_27_<5>) );
	DFFPOSX1 DFFPOSX1_615 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3676), .Q(dp.rf.rf_27_<6>) );
	DFFPOSX1 DFFPOSX1_616 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3677), .Q(dp.rf.rf_27_<7>) );
	DFFPOSX1 DFFPOSX1_617 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3678), .Q(dp.rf.rf_27_<8>) );
	DFFPOSX1 DFFPOSX1_618 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3679), .Q(dp.rf.rf_27_<9>) );
	DFFPOSX1 DFFPOSX1_619 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3680), .Q(dp.rf.rf_27_<10>) );
	DFFPOSX1 DFFPOSX1_620 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3681), .Q(dp.rf.rf_27_<11>) );
	DFFPOSX1 DFFPOSX1_621 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3682), .Q(dp.rf.rf_27_<12>) );
	DFFPOSX1 DFFPOSX1_622 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3683), .Q(dp.rf.rf_27_<13>) );
	DFFPOSX1 DFFPOSX1_623 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3684), .Q(dp.rf.rf_27_<14>) );
	DFFPOSX1 DFFPOSX1_624 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3685), .Q(dp.rf.rf_27_<15>) );
	DFFPOSX1 DFFPOSX1_625 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3686), .Q(dp.rf.rf_27_<16>) );
	DFFPOSX1 DFFPOSX1_626 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3687), .Q(dp.rf.rf_27_<17>) );
	DFFPOSX1 DFFPOSX1_627 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3688), .Q(dp.rf.rf_27_<18>) );
	DFFPOSX1 DFFPOSX1_628 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3689), .Q(dp.rf.rf_27_<19>) );
	DFFPOSX1 DFFPOSX1_629 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3690), .Q(dp.rf.rf_27_<20>) );
	DFFPOSX1 DFFPOSX1_630 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3691), .Q(dp.rf.rf_27_<21>) );
	DFFPOSX1 DFFPOSX1_631 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3692), .Q(dp.rf.rf_27_<22>) );
	DFFPOSX1 DFFPOSX1_632 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3693), .Q(dp.rf.rf_27_<23>) );
	DFFPOSX1 DFFPOSX1_633 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3694), .Q(dp.rf.rf_27_<24>) );
	DFFPOSX1 DFFPOSX1_634 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3695), .Q(dp.rf.rf_27_<25>) );
	DFFPOSX1 DFFPOSX1_635 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3696), .Q(dp.rf.rf_27_<26>) );
	DFFPOSX1 DFFPOSX1_636 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3697), .Q(dp.rf.rf_27_<27>) );
	DFFPOSX1 DFFPOSX1_637 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3698), .Q(dp.rf.rf_27_<28>) );
	DFFPOSX1 DFFPOSX1_638 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3699), .Q(dp.rf.rf_27_<29>) );
	DFFPOSX1 DFFPOSX1_639 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3700), .Q(dp.rf.rf_27_<30>) );
	DFFPOSX1 DFFPOSX1_640 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3701), .Q(dp.rf.rf_27_<31>) );
	DFFPOSX1 DFFPOSX1_641 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3702), .Q(dp.rf.rf_28_<0>) );
	DFFPOSX1 DFFPOSX1_642 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3703), .Q(dp.rf.rf_28_<1>) );
	DFFPOSX1 DFFPOSX1_643 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3704), .Q(dp.rf.rf_28_<2>) );
	DFFPOSX1 DFFPOSX1_644 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3705), .Q(dp.rf.rf_28_<3>) );
	DFFPOSX1 DFFPOSX1_645 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3706), .Q(dp.rf.rf_28_<4>) );
	DFFPOSX1 DFFPOSX1_646 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3707), .Q(dp.rf.rf_28_<5>) );
	DFFPOSX1 DFFPOSX1_647 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3708), .Q(dp.rf.rf_28_<6>) );
	DFFPOSX1 DFFPOSX1_648 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3709), .Q(dp.rf.rf_28_<7>) );
	DFFPOSX1 DFFPOSX1_649 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3710), .Q(dp.rf.rf_28_<8>) );
	DFFPOSX1 DFFPOSX1_650 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3711), .Q(dp.rf.rf_28_<9>) );
	DFFPOSX1 DFFPOSX1_651 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3712), .Q(dp.rf.rf_28_<10>) );
	DFFPOSX1 DFFPOSX1_652 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3713), .Q(dp.rf.rf_28_<11>) );
	DFFPOSX1 DFFPOSX1_653 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3714), .Q(dp.rf.rf_28_<12>) );
	DFFPOSX1 DFFPOSX1_654 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3715), .Q(dp.rf.rf_28_<13>) );
	DFFPOSX1 DFFPOSX1_655 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3716), .Q(dp.rf.rf_28_<14>) );
	DFFPOSX1 DFFPOSX1_656 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3717), .Q(dp.rf.rf_28_<15>) );
	DFFPOSX1 DFFPOSX1_657 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3718), .Q(dp.rf.rf_28_<16>) );
	DFFPOSX1 DFFPOSX1_658 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3719), .Q(dp.rf.rf_28_<17>) );
	DFFPOSX1 DFFPOSX1_659 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3720), .Q(dp.rf.rf_28_<18>) );
	DFFPOSX1 DFFPOSX1_660 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3721), .Q(dp.rf.rf_28_<19>) );
	DFFPOSX1 DFFPOSX1_661 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3722), .Q(dp.rf.rf_28_<20>) );
	DFFPOSX1 DFFPOSX1_662 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3723), .Q(dp.rf.rf_28_<21>) );
	DFFPOSX1 DFFPOSX1_663 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3724), .Q(dp.rf.rf_28_<22>) );
	DFFPOSX1 DFFPOSX1_664 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3725), .Q(dp.rf.rf_28_<23>) );
	DFFPOSX1 DFFPOSX1_665 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3726), .Q(dp.rf.rf_28_<24>) );
	DFFPOSX1 DFFPOSX1_666 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3727), .Q(dp.rf.rf_28_<25>) );
	DFFPOSX1 DFFPOSX1_667 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3728), .Q(dp.rf.rf_28_<26>) );
	DFFPOSX1 DFFPOSX1_668 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3729), .Q(dp.rf.rf_28_<27>) );
	DFFPOSX1 DFFPOSX1_669 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3730), .Q(dp.rf.rf_28_<28>) );
	DFFPOSX1 DFFPOSX1_670 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3731), .Q(dp.rf.rf_28_<29>) );
	DFFPOSX1 DFFPOSX1_671 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3732), .Q(dp.rf.rf_28_<30>) );
	DFFPOSX1 DFFPOSX1_672 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3733), .Q(dp.rf.rf_28_<31>) );
	DFFPOSX1 DFFPOSX1_673 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3734), .Q(dp.rf.rf_29_<0>) );
	DFFPOSX1 DFFPOSX1_674 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3735), .Q(dp.rf.rf_29_<1>) );
	DFFPOSX1 DFFPOSX1_675 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3736), .Q(dp.rf.rf_29_<2>) );
	DFFPOSX1 DFFPOSX1_676 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3737), .Q(dp.rf.rf_29_<3>) );
	DFFPOSX1 DFFPOSX1_677 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3738), .Q(dp.rf.rf_29_<4>) );
	DFFPOSX1 DFFPOSX1_678 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3739), .Q(dp.rf.rf_29_<5>) );
	DFFPOSX1 DFFPOSX1_679 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3740), .Q(dp.rf.rf_29_<6>) );
	DFFPOSX1 DFFPOSX1_680 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3741), .Q(dp.rf.rf_29_<7>) );
	DFFPOSX1 DFFPOSX1_681 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3742), .Q(dp.rf.rf_29_<8>) );
	DFFPOSX1 DFFPOSX1_682 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3743), .Q(dp.rf.rf_29_<9>) );
	DFFPOSX1 DFFPOSX1_683 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3744), .Q(dp.rf.rf_29_<10>) );
	DFFPOSX1 DFFPOSX1_684 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3745), .Q(dp.rf.rf_29_<11>) );
	DFFPOSX1 DFFPOSX1_685 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3746), .Q(dp.rf.rf_29_<12>) );
	DFFPOSX1 DFFPOSX1_686 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3747), .Q(dp.rf.rf_29_<13>) );
	DFFPOSX1 DFFPOSX1_687 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3748), .Q(dp.rf.rf_29_<14>) );
	DFFPOSX1 DFFPOSX1_688 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3749), .Q(dp.rf.rf_29_<15>) );
	DFFPOSX1 DFFPOSX1_689 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3750), .Q(dp.rf.rf_29_<16>) );
	DFFPOSX1 DFFPOSX1_690 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3751), .Q(dp.rf.rf_29_<17>) );
	DFFPOSX1 DFFPOSX1_691 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3752), .Q(dp.rf.rf_29_<18>) );
	DFFPOSX1 DFFPOSX1_692 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3753), .Q(dp.rf.rf_29_<19>) );
	DFFPOSX1 DFFPOSX1_693 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3754), .Q(dp.rf.rf_29_<20>) );
	DFFPOSX1 DFFPOSX1_694 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3755), .Q(dp.rf.rf_29_<21>) );
	DFFPOSX1 DFFPOSX1_695 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3756), .Q(dp.rf.rf_29_<22>) );
	DFFPOSX1 DFFPOSX1_696 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3757), .Q(dp.rf.rf_29_<23>) );
	DFFPOSX1 DFFPOSX1_697 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3758), .Q(dp.rf.rf_29_<24>) );
	DFFPOSX1 DFFPOSX1_698 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3759), .Q(dp.rf.rf_29_<25>) );
	DFFPOSX1 DFFPOSX1_699 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3760), .Q(dp.rf.rf_29_<26>) );
	DFFPOSX1 DFFPOSX1_700 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3761), .Q(dp.rf.rf_29_<27>) );
	DFFPOSX1 DFFPOSX1_701 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3762), .Q(dp.rf.rf_29_<28>) );
	DFFPOSX1 DFFPOSX1_702 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3763), .Q(dp.rf.rf_29_<29>) );
	DFFPOSX1 DFFPOSX1_703 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3764), .Q(dp.rf.rf_29_<30>) );
	DFFPOSX1 DFFPOSX1_704 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3765), .Q(dp.rf.rf_29_<31>) );
	DFFPOSX1 DFFPOSX1_705 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3766), .Q(dp.rf.rf_2_<0>) );
	DFFPOSX1 DFFPOSX1_706 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3767), .Q(dp.rf.rf_2_<1>) );
	DFFPOSX1 DFFPOSX1_707 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3768), .Q(dp.rf.rf_2_<2>) );
	DFFPOSX1 DFFPOSX1_708 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3769), .Q(dp.rf.rf_2_<3>) );
	DFFPOSX1 DFFPOSX1_709 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3770), .Q(dp.rf.rf_2_<4>) );
	DFFPOSX1 DFFPOSX1_710 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3771), .Q(dp.rf.rf_2_<5>) );
	DFFPOSX1 DFFPOSX1_711 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3772), .Q(dp.rf.rf_2_<6>) );
	DFFPOSX1 DFFPOSX1_712 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3773), .Q(dp.rf.rf_2_<7>) );
	DFFPOSX1 DFFPOSX1_713 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3774), .Q(dp.rf.rf_2_<8>) );
	DFFPOSX1 DFFPOSX1_714 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3775), .Q(dp.rf.rf_2_<9>) );
	DFFPOSX1 DFFPOSX1_715 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3776), .Q(dp.rf.rf_2_<10>) );
	DFFPOSX1 DFFPOSX1_716 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3777), .Q(dp.rf.rf_2_<11>) );
	DFFPOSX1 DFFPOSX1_717 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3778), .Q(dp.rf.rf_2_<12>) );
	DFFPOSX1 DFFPOSX1_718 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3779), .Q(dp.rf.rf_2_<13>) );
	DFFPOSX1 DFFPOSX1_719 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3780), .Q(dp.rf.rf_2_<14>) );
	DFFPOSX1 DFFPOSX1_720 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3781), .Q(dp.rf.rf_2_<15>) );
	DFFPOSX1 DFFPOSX1_721 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3782), .Q(dp.rf.rf_2_<16>) );
	DFFPOSX1 DFFPOSX1_722 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3783), .Q(dp.rf.rf_2_<17>) );
	DFFPOSX1 DFFPOSX1_723 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3784), .Q(dp.rf.rf_2_<18>) );
	DFFPOSX1 DFFPOSX1_724 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3785), .Q(dp.rf.rf_2_<19>) );
	DFFPOSX1 DFFPOSX1_725 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3786), .Q(dp.rf.rf_2_<20>) );
	DFFPOSX1 DFFPOSX1_726 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3787), .Q(dp.rf.rf_2_<21>) );
	DFFPOSX1 DFFPOSX1_727 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3788), .Q(dp.rf.rf_2_<22>) );
	DFFPOSX1 DFFPOSX1_728 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3789), .Q(dp.rf.rf_2_<23>) );
	DFFPOSX1 DFFPOSX1_729 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3790), .Q(dp.rf.rf_2_<24>) );
	DFFPOSX1 DFFPOSX1_730 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3791), .Q(dp.rf.rf_2_<25>) );
	DFFPOSX1 DFFPOSX1_731 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3792), .Q(dp.rf.rf_2_<26>) );
	DFFPOSX1 DFFPOSX1_732 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3793), .Q(dp.rf.rf_2_<27>) );
	DFFPOSX1 DFFPOSX1_733 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3794), .Q(dp.rf.rf_2_<28>) );
	DFFPOSX1 DFFPOSX1_734 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3795), .Q(dp.rf.rf_2_<29>) );
	DFFPOSX1 DFFPOSX1_735 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3796), .Q(dp.rf.rf_2_<30>) );
	DFFPOSX1 DFFPOSX1_736 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3797), .Q(dp.rf.rf_2_<31>) );
	DFFPOSX1 DFFPOSX1_737 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3798), .Q(dp.rf.rf_30_<0>) );
	DFFPOSX1 DFFPOSX1_738 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3799), .Q(dp.rf.rf_30_<1>) );
	DFFPOSX1 DFFPOSX1_739 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3800), .Q(dp.rf.rf_30_<2>) );
	DFFPOSX1 DFFPOSX1_740 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3801), .Q(dp.rf.rf_30_<3>) );
	DFFPOSX1 DFFPOSX1_741 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3802), .Q(dp.rf.rf_30_<4>) );
	DFFPOSX1 DFFPOSX1_742 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3803), .Q(dp.rf.rf_30_<5>) );
	DFFPOSX1 DFFPOSX1_743 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3804), .Q(dp.rf.rf_30_<6>) );
	DFFPOSX1 DFFPOSX1_744 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3805), .Q(dp.rf.rf_30_<7>) );
	DFFPOSX1 DFFPOSX1_745 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3806), .Q(dp.rf.rf_30_<8>) );
	DFFPOSX1 DFFPOSX1_746 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3807), .Q(dp.rf.rf_30_<9>) );
	DFFPOSX1 DFFPOSX1_747 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3808), .Q(dp.rf.rf_30_<10>) );
	DFFPOSX1 DFFPOSX1_748 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3809), .Q(dp.rf.rf_30_<11>) );
	DFFPOSX1 DFFPOSX1_749 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3810), .Q(dp.rf.rf_30_<12>) );
	DFFPOSX1 DFFPOSX1_750 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3811), .Q(dp.rf.rf_30_<13>) );
	DFFPOSX1 DFFPOSX1_751 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3812), .Q(dp.rf.rf_30_<14>) );
	DFFPOSX1 DFFPOSX1_752 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3813), .Q(dp.rf.rf_30_<15>) );
	DFFPOSX1 DFFPOSX1_753 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3814), .Q(dp.rf.rf_30_<16>) );
	DFFPOSX1 DFFPOSX1_754 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3815), .Q(dp.rf.rf_30_<17>) );
	DFFPOSX1 DFFPOSX1_755 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3816), .Q(dp.rf.rf_30_<18>) );
	DFFPOSX1 DFFPOSX1_756 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3817), .Q(dp.rf.rf_30_<19>) );
	DFFPOSX1 DFFPOSX1_757 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3818), .Q(dp.rf.rf_30_<20>) );
	DFFPOSX1 DFFPOSX1_758 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3819), .Q(dp.rf.rf_30_<21>) );
	DFFPOSX1 DFFPOSX1_759 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3820), .Q(dp.rf.rf_30_<22>) );
	DFFPOSX1 DFFPOSX1_760 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3821), .Q(dp.rf.rf_30_<23>) );
	DFFPOSX1 DFFPOSX1_761 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3822), .Q(dp.rf.rf_30_<24>) );
	DFFPOSX1 DFFPOSX1_762 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3823), .Q(dp.rf.rf_30_<25>) );
	DFFPOSX1 DFFPOSX1_763 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3824), .Q(dp.rf.rf_30_<26>) );
	DFFPOSX1 DFFPOSX1_764 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3825), .Q(dp.rf.rf_30_<27>) );
	DFFPOSX1 DFFPOSX1_765 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3826), .Q(dp.rf.rf_30_<28>) );
	DFFPOSX1 DFFPOSX1_766 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3827), .Q(dp.rf.rf_30_<29>) );
	DFFPOSX1 DFFPOSX1_767 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3828), .Q(dp.rf.rf_30_<30>) );
	DFFPOSX1 DFFPOSX1_768 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3829), .Q(dp.rf.rf_30_<31>) );
	DFFPOSX1 DFFPOSX1_769 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3830), .Q(dp.rf.rf_31_<0>) );
	DFFPOSX1 DFFPOSX1_770 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3831), .Q(dp.rf.rf_31_<1>) );
	DFFPOSX1 DFFPOSX1_771 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3832), .Q(dp.rf.rf_31_<2>) );
	DFFPOSX1 DFFPOSX1_772 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3833), .Q(dp.rf.rf_31_<3>) );
	DFFPOSX1 DFFPOSX1_773 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3834), .Q(dp.rf.rf_31_<4>) );
	DFFPOSX1 DFFPOSX1_774 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3835), .Q(dp.rf.rf_31_<5>) );
	DFFPOSX1 DFFPOSX1_775 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3836), .Q(dp.rf.rf_31_<6>) );
	DFFPOSX1 DFFPOSX1_776 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3837), .Q(dp.rf.rf_31_<7>) );
	DFFPOSX1 DFFPOSX1_777 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3838), .Q(dp.rf.rf_31_<8>) );
	DFFPOSX1 DFFPOSX1_778 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3839), .Q(dp.rf.rf_31_<9>) );
	DFFPOSX1 DFFPOSX1_779 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3840), .Q(dp.rf.rf_31_<10>) );
	DFFPOSX1 DFFPOSX1_780 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3841), .Q(dp.rf.rf_31_<11>) );
	DFFPOSX1 DFFPOSX1_781 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3842), .Q(dp.rf.rf_31_<12>) );
	DFFPOSX1 DFFPOSX1_782 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3843), .Q(dp.rf.rf_31_<13>) );
	DFFPOSX1 DFFPOSX1_783 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3844), .Q(dp.rf.rf_31_<14>) );
	DFFPOSX1 DFFPOSX1_784 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3845), .Q(dp.rf.rf_31_<15>) );
	DFFPOSX1 DFFPOSX1_785 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3846), .Q(dp.rf.rf_31_<16>) );
	DFFPOSX1 DFFPOSX1_786 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3847), .Q(dp.rf.rf_31_<17>) );
	DFFPOSX1 DFFPOSX1_787 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3848), .Q(dp.rf.rf_31_<18>) );
	DFFPOSX1 DFFPOSX1_788 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3849), .Q(dp.rf.rf_31_<19>) );
	DFFPOSX1 DFFPOSX1_789 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3850), .Q(dp.rf.rf_31_<20>) );
	DFFPOSX1 DFFPOSX1_790 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3851), .Q(dp.rf.rf_31_<21>) );
	DFFPOSX1 DFFPOSX1_791 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3852), .Q(dp.rf.rf_31_<22>) );
	DFFPOSX1 DFFPOSX1_792 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3853), .Q(dp.rf.rf_31_<23>) );
	DFFPOSX1 DFFPOSX1_793 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3854), .Q(dp.rf.rf_31_<24>) );
	DFFPOSX1 DFFPOSX1_794 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3855), .Q(dp.rf.rf_31_<25>) );
	DFFPOSX1 DFFPOSX1_795 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3856), .Q(dp.rf.rf_31_<26>) );
	DFFPOSX1 DFFPOSX1_796 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3857), .Q(dp.rf.rf_31_<27>) );
	DFFPOSX1 DFFPOSX1_797 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3858), .Q(dp.rf.rf_31_<28>) );
	DFFPOSX1 DFFPOSX1_798 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3859), .Q(dp.rf.rf_31_<29>) );
	DFFPOSX1 DFFPOSX1_799 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3860), .Q(dp.rf.rf_31_<30>) );
	DFFPOSX1 DFFPOSX1_800 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3861), .Q(dp.rf.rf_31_<31>) );
	DFFPOSX1 DFFPOSX1_801 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3862), .Q(dp.rf.rf_3_<0>) );
	DFFPOSX1 DFFPOSX1_802 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3863), .Q(dp.rf.rf_3_<1>) );
	DFFPOSX1 DFFPOSX1_803 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3864), .Q(dp.rf.rf_3_<2>) );
	DFFPOSX1 DFFPOSX1_804 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3865), .Q(dp.rf.rf_3_<3>) );
	DFFPOSX1 DFFPOSX1_805 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3866), .Q(dp.rf.rf_3_<4>) );
	DFFPOSX1 DFFPOSX1_806 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3867), .Q(dp.rf.rf_3_<5>) );
	DFFPOSX1 DFFPOSX1_807 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3868), .Q(dp.rf.rf_3_<6>) );
	DFFPOSX1 DFFPOSX1_808 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3869), .Q(dp.rf.rf_3_<7>) );
	DFFPOSX1 DFFPOSX1_809 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3870), .Q(dp.rf.rf_3_<8>) );
	DFFPOSX1 DFFPOSX1_810 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3871), .Q(dp.rf.rf_3_<9>) );
	DFFPOSX1 DFFPOSX1_811 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3872), .Q(dp.rf.rf_3_<10>) );
	DFFPOSX1 DFFPOSX1_812 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3873), .Q(dp.rf.rf_3_<11>) );
	DFFPOSX1 DFFPOSX1_813 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3874), .Q(dp.rf.rf_3_<12>) );
	DFFPOSX1 DFFPOSX1_814 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3875), .Q(dp.rf.rf_3_<13>) );
	DFFPOSX1 DFFPOSX1_815 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3876), .Q(dp.rf.rf_3_<14>) );
	DFFPOSX1 DFFPOSX1_816 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3877), .Q(dp.rf.rf_3_<15>) );
	DFFPOSX1 DFFPOSX1_817 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3878), .Q(dp.rf.rf_3_<16>) );
	DFFPOSX1 DFFPOSX1_818 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3879), .Q(dp.rf.rf_3_<17>) );
	DFFPOSX1 DFFPOSX1_819 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3880), .Q(dp.rf.rf_3_<18>) );
	DFFPOSX1 DFFPOSX1_820 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3881), .Q(dp.rf.rf_3_<19>) );
	DFFPOSX1 DFFPOSX1_821 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3882), .Q(dp.rf.rf_3_<20>) );
	DFFPOSX1 DFFPOSX1_822 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3883), .Q(dp.rf.rf_3_<21>) );
	DFFPOSX1 DFFPOSX1_823 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3884), .Q(dp.rf.rf_3_<22>) );
	DFFPOSX1 DFFPOSX1_824 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3885), .Q(dp.rf.rf_3_<23>) );
	DFFPOSX1 DFFPOSX1_825 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3886), .Q(dp.rf.rf_3_<24>) );
	DFFPOSX1 DFFPOSX1_826 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3887), .Q(dp.rf.rf_3_<25>) );
	DFFPOSX1 DFFPOSX1_827 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3888), .Q(dp.rf.rf_3_<26>) );
	DFFPOSX1 DFFPOSX1_828 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3889), .Q(dp.rf.rf_3_<27>) );
	DFFPOSX1 DFFPOSX1_829 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3890), .Q(dp.rf.rf_3_<28>) );
	DFFPOSX1 DFFPOSX1_830 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3891), .Q(dp.rf.rf_3_<29>) );
	DFFPOSX1 DFFPOSX1_831 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3892), .Q(dp.rf.rf_3_<30>) );
	DFFPOSX1 DFFPOSX1_832 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3893), .Q(dp.rf.rf_3_<31>) );
	DFFPOSX1 DFFPOSX1_833 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3894), .Q(dp.rf.rf_4_<0>) );
	DFFPOSX1 DFFPOSX1_834 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3895), .Q(dp.rf.rf_4_<1>) );
	DFFPOSX1 DFFPOSX1_835 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3896), .Q(dp.rf.rf_4_<2>) );
	DFFPOSX1 DFFPOSX1_836 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3897), .Q(dp.rf.rf_4_<3>) );
	DFFPOSX1 DFFPOSX1_837 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3898), .Q(dp.rf.rf_4_<4>) );
	DFFPOSX1 DFFPOSX1_838 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3899), .Q(dp.rf.rf_4_<5>) );
	DFFPOSX1 DFFPOSX1_839 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3900), .Q(dp.rf.rf_4_<6>) );
	DFFPOSX1 DFFPOSX1_840 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3901), .Q(dp.rf.rf_4_<7>) );
	DFFPOSX1 DFFPOSX1_841 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3902), .Q(dp.rf.rf_4_<8>) );
	DFFPOSX1 DFFPOSX1_842 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3903), .Q(dp.rf.rf_4_<9>) );
	DFFPOSX1 DFFPOSX1_843 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3904), .Q(dp.rf.rf_4_<10>) );
	DFFPOSX1 DFFPOSX1_844 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3905), .Q(dp.rf.rf_4_<11>) );
	DFFPOSX1 DFFPOSX1_845 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3906), .Q(dp.rf.rf_4_<12>) );
	DFFPOSX1 DFFPOSX1_846 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3907), .Q(dp.rf.rf_4_<13>) );
	DFFPOSX1 DFFPOSX1_847 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3908), .Q(dp.rf.rf_4_<14>) );
	DFFPOSX1 DFFPOSX1_848 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3909), .Q(dp.rf.rf_4_<15>) );
	DFFPOSX1 DFFPOSX1_849 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3910), .Q(dp.rf.rf_4_<16>) );
	DFFPOSX1 DFFPOSX1_850 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3911), .Q(dp.rf.rf_4_<17>) );
	DFFPOSX1 DFFPOSX1_851 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3912), .Q(dp.rf.rf_4_<18>) );
	DFFPOSX1 DFFPOSX1_852 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3913), .Q(dp.rf.rf_4_<19>) );
	DFFPOSX1 DFFPOSX1_853 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3914), .Q(dp.rf.rf_4_<20>) );
	DFFPOSX1 DFFPOSX1_854 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3915), .Q(dp.rf.rf_4_<21>) );
	DFFPOSX1 DFFPOSX1_855 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3916), .Q(dp.rf.rf_4_<22>) );
	DFFPOSX1 DFFPOSX1_856 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3917), .Q(dp.rf.rf_4_<23>) );
	DFFPOSX1 DFFPOSX1_857 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3918), .Q(dp.rf.rf_4_<24>) );
	DFFPOSX1 DFFPOSX1_858 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3919), .Q(dp.rf.rf_4_<25>) );
	DFFPOSX1 DFFPOSX1_859 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3920), .Q(dp.rf.rf_4_<26>) );
	DFFPOSX1 DFFPOSX1_860 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3921), .Q(dp.rf.rf_4_<27>) );
	DFFPOSX1 DFFPOSX1_861 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3922), .Q(dp.rf.rf_4_<28>) );
	DFFPOSX1 DFFPOSX1_862 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3923), .Q(dp.rf.rf_4_<29>) );
	DFFPOSX1 DFFPOSX1_863 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3924), .Q(dp.rf.rf_4_<30>) );
	DFFPOSX1 DFFPOSX1_864 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3925), .Q(dp.rf.rf_4_<31>) );
	DFFPOSX1 DFFPOSX1_865 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3926), .Q(dp.rf.rf_5_<0>) );
	DFFPOSX1 DFFPOSX1_866 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3927), .Q(dp.rf.rf_5_<1>) );
	DFFPOSX1 DFFPOSX1_867 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3928), .Q(dp.rf.rf_5_<2>) );
	DFFPOSX1 DFFPOSX1_868 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3929), .Q(dp.rf.rf_5_<3>) );
	DFFPOSX1 DFFPOSX1_869 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3930), .Q(dp.rf.rf_5_<4>) );
	DFFPOSX1 DFFPOSX1_870 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3931), .Q(dp.rf.rf_5_<5>) );
	DFFPOSX1 DFFPOSX1_871 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3932), .Q(dp.rf.rf_5_<6>) );
	DFFPOSX1 DFFPOSX1_872 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3933), .Q(dp.rf.rf_5_<7>) );
	DFFPOSX1 DFFPOSX1_873 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3934), .Q(dp.rf.rf_5_<8>) );
	DFFPOSX1 DFFPOSX1_874 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3935), .Q(dp.rf.rf_5_<9>) );
	DFFPOSX1 DFFPOSX1_875 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3936), .Q(dp.rf.rf_5_<10>) );
	DFFPOSX1 DFFPOSX1_876 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3937), .Q(dp.rf.rf_5_<11>) );
	DFFPOSX1 DFFPOSX1_877 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3938), .Q(dp.rf.rf_5_<12>) );
	DFFPOSX1 DFFPOSX1_878 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3939), .Q(dp.rf.rf_5_<13>) );
	DFFPOSX1 DFFPOSX1_879 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3940), .Q(dp.rf.rf_5_<14>) );
	DFFPOSX1 DFFPOSX1_880 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3941), .Q(dp.rf.rf_5_<15>) );
	DFFPOSX1 DFFPOSX1_881 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3942), .Q(dp.rf.rf_5_<16>) );
	DFFPOSX1 DFFPOSX1_882 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3943), .Q(dp.rf.rf_5_<17>) );
	DFFPOSX1 DFFPOSX1_883 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3944), .Q(dp.rf.rf_5_<18>) );
	DFFPOSX1 DFFPOSX1_884 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3945), .Q(dp.rf.rf_5_<19>) );
	DFFPOSX1 DFFPOSX1_885 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3946), .Q(dp.rf.rf_5_<20>) );
	DFFPOSX1 DFFPOSX1_886 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3947), .Q(dp.rf.rf_5_<21>) );
	DFFPOSX1 DFFPOSX1_887 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3948), .Q(dp.rf.rf_5_<22>) );
	DFFPOSX1 DFFPOSX1_888 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3949), .Q(dp.rf.rf_5_<23>) );
	DFFPOSX1 DFFPOSX1_889 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3950), .Q(dp.rf.rf_5_<24>) );
	DFFPOSX1 DFFPOSX1_890 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3951), .Q(dp.rf.rf_5_<25>) );
	DFFPOSX1 DFFPOSX1_891 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3952), .Q(dp.rf.rf_5_<26>) );
	DFFPOSX1 DFFPOSX1_892 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3953), .Q(dp.rf.rf_5_<27>) );
	DFFPOSX1 DFFPOSX1_893 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3954), .Q(dp.rf.rf_5_<28>) );
	DFFPOSX1 DFFPOSX1_894 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3955), .Q(dp.rf.rf_5_<29>) );
	DFFPOSX1 DFFPOSX1_895 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3956), .Q(dp.rf.rf_5_<30>) );
	DFFPOSX1 DFFPOSX1_896 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3957), .Q(dp.rf.rf_5_<31>) );
	DFFPOSX1 DFFPOSX1_897 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3958), .Q(dp.rf.rf_6_<0>) );
	DFFPOSX1 DFFPOSX1_898 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3959), .Q(dp.rf.rf_6_<1>) );
	DFFPOSX1 DFFPOSX1_899 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3960), .Q(dp.rf.rf_6_<2>) );
	DFFPOSX1 DFFPOSX1_900 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3961), .Q(dp.rf.rf_6_<3>) );
	DFFPOSX1 DFFPOSX1_901 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3962), .Q(dp.rf.rf_6_<4>) );
	DFFPOSX1 DFFPOSX1_902 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3963), .Q(dp.rf.rf_6_<5>) );
	DFFPOSX1 DFFPOSX1_903 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3964), .Q(dp.rf.rf_6_<6>) );
	DFFPOSX1 DFFPOSX1_904 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3965), .Q(dp.rf.rf_6_<7>) );
	DFFPOSX1 DFFPOSX1_905 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3966), .Q(dp.rf.rf_6_<8>) );
	DFFPOSX1 DFFPOSX1_906 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3967), .Q(dp.rf.rf_6_<9>) );
	DFFPOSX1 DFFPOSX1_907 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3968), .Q(dp.rf.rf_6_<10>) );
	DFFPOSX1 DFFPOSX1_908 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3969), .Q(dp.rf.rf_6_<11>) );
	DFFPOSX1 DFFPOSX1_909 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3970), .Q(dp.rf.rf_6_<12>) );
	DFFPOSX1 DFFPOSX1_910 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3971), .Q(dp.rf.rf_6_<13>) );
	DFFPOSX1 DFFPOSX1_911 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3972), .Q(dp.rf.rf_6_<14>) );
	DFFPOSX1 DFFPOSX1_912 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3973), .Q(dp.rf.rf_6_<15>) );
	DFFPOSX1 DFFPOSX1_913 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3974), .Q(dp.rf.rf_6_<16>) );
	DFFPOSX1 DFFPOSX1_914 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3975), .Q(dp.rf.rf_6_<17>) );
	DFFPOSX1 DFFPOSX1_915 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3976), .Q(dp.rf.rf_6_<18>) );
	DFFPOSX1 DFFPOSX1_916 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3977), .Q(dp.rf.rf_6_<19>) );
	DFFPOSX1 DFFPOSX1_917 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3978), .Q(dp.rf.rf_6_<20>) );
	DFFPOSX1 DFFPOSX1_918 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3979), .Q(dp.rf.rf_6_<21>) );
	DFFPOSX1 DFFPOSX1_919 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3980), .Q(dp.rf.rf_6_<22>) );
	DFFPOSX1 DFFPOSX1_920 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3981), .Q(dp.rf.rf_6_<23>) );
	DFFPOSX1 DFFPOSX1_921 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3982), .Q(dp.rf.rf_6_<24>) );
	DFFPOSX1 DFFPOSX1_922 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3983), .Q(dp.rf.rf_6_<25>) );
	DFFPOSX1 DFFPOSX1_923 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3984), .Q(dp.rf.rf_6_<26>) );
	DFFPOSX1 DFFPOSX1_924 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3985), .Q(dp.rf.rf_6_<27>) );
	DFFPOSX1 DFFPOSX1_925 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3986), .Q(dp.rf.rf_6_<28>) );
	DFFPOSX1 DFFPOSX1_926 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3987), .Q(dp.rf.rf_6_<29>) );
	DFFPOSX1 DFFPOSX1_927 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3988), .Q(dp.rf.rf_6_<30>) );
	DFFPOSX1 DFFPOSX1_928 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3989), .Q(dp.rf.rf_6_<31>) );
	DFFPOSX1 DFFPOSX1_929 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3990), .Q(dp.rf.rf_7_<0>) );
	DFFPOSX1 DFFPOSX1_930 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3991), .Q(dp.rf.rf_7_<1>) );
	DFFPOSX1 DFFPOSX1_931 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3992), .Q(dp.rf.rf_7_<2>) );
	DFFPOSX1 DFFPOSX1_932 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3993), .Q(dp.rf.rf_7_<3>) );
	DFFPOSX1 DFFPOSX1_933 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3994), .Q(dp.rf.rf_7_<4>) );
	DFFPOSX1 DFFPOSX1_934 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3995), .Q(dp.rf.rf_7_<5>) );
	DFFPOSX1 DFFPOSX1_935 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3996), .Q(dp.rf.rf_7_<6>) );
	DFFPOSX1 DFFPOSX1_936 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3997), .Q(dp.rf.rf_7_<7>) );
	DFFPOSX1 DFFPOSX1_937 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3998), .Q(dp.rf.rf_7_<8>) );
	DFFPOSX1 DFFPOSX1_938 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n3999), .Q(dp.rf.rf_7_<9>) );
	DFFPOSX1 DFFPOSX1_939 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4000), .Q(dp.rf.rf_7_<10>) );
	DFFPOSX1 DFFPOSX1_940 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4001), .Q(dp.rf.rf_7_<11>) );
	DFFPOSX1 DFFPOSX1_941 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4002), .Q(dp.rf.rf_7_<12>) );
	DFFPOSX1 DFFPOSX1_942 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4003), .Q(dp.rf.rf_7_<13>) );
	DFFPOSX1 DFFPOSX1_943 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4004), .Q(dp.rf.rf_7_<14>) );
	DFFPOSX1 DFFPOSX1_944 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4005), .Q(dp.rf.rf_7_<15>) );
	DFFPOSX1 DFFPOSX1_945 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4006), .Q(dp.rf.rf_7_<16>) );
	DFFPOSX1 DFFPOSX1_946 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4007), .Q(dp.rf.rf_7_<17>) );
	DFFPOSX1 DFFPOSX1_947 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4008), .Q(dp.rf.rf_7_<18>) );
	DFFPOSX1 DFFPOSX1_948 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4009), .Q(dp.rf.rf_7_<19>) );
	DFFPOSX1 DFFPOSX1_949 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4010), .Q(dp.rf.rf_7_<20>) );
	DFFPOSX1 DFFPOSX1_950 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4011), .Q(dp.rf.rf_7_<21>) );
	DFFPOSX1 DFFPOSX1_951 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4012), .Q(dp.rf.rf_7_<22>) );
	DFFPOSX1 DFFPOSX1_952 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4013), .Q(dp.rf.rf_7_<23>) );
	DFFPOSX1 DFFPOSX1_953 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4014), .Q(dp.rf.rf_7_<24>) );
	DFFPOSX1 DFFPOSX1_954 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4015), .Q(dp.rf.rf_7_<25>) );
	DFFPOSX1 DFFPOSX1_955 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4016), .Q(dp.rf.rf_7_<26>) );
	DFFPOSX1 DFFPOSX1_956 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4017), .Q(dp.rf.rf_7_<27>) );
	DFFPOSX1 DFFPOSX1_957 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4018), .Q(dp.rf.rf_7_<28>) );
	DFFPOSX1 DFFPOSX1_958 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4019), .Q(dp.rf.rf_7_<29>) );
	DFFPOSX1 DFFPOSX1_959 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4020), .Q(dp.rf.rf_7_<30>) );
	DFFPOSX1 DFFPOSX1_960 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4021), .Q(dp.rf.rf_7_<31>) );
	DFFPOSX1 DFFPOSX1_961 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4022), .Q(dp.rf.rf_8_<0>) );
	DFFPOSX1 DFFPOSX1_962 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4023), .Q(dp.rf.rf_8_<1>) );
	DFFPOSX1 DFFPOSX1_963 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4024), .Q(dp.rf.rf_8_<2>) );
	DFFPOSX1 DFFPOSX1_964 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4025), .Q(dp.rf.rf_8_<3>) );
	DFFPOSX1 DFFPOSX1_965 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4026), .Q(dp.rf.rf_8_<4>) );
	DFFPOSX1 DFFPOSX1_966 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4027), .Q(dp.rf.rf_8_<5>) );
	DFFPOSX1 DFFPOSX1_967 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4028), .Q(dp.rf.rf_8_<6>) );
	DFFPOSX1 DFFPOSX1_968 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4029), .Q(dp.rf.rf_8_<7>) );
	DFFPOSX1 DFFPOSX1_969 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4030), .Q(dp.rf.rf_8_<8>) );
	DFFPOSX1 DFFPOSX1_970 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4031), .Q(dp.rf.rf_8_<9>) );
	DFFPOSX1 DFFPOSX1_971 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4032), .Q(dp.rf.rf_8_<10>) );
	DFFPOSX1 DFFPOSX1_972 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4033), .Q(dp.rf.rf_8_<11>) );
	DFFPOSX1 DFFPOSX1_973 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4034), .Q(dp.rf.rf_8_<12>) );
	DFFPOSX1 DFFPOSX1_974 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4035), .Q(dp.rf.rf_8_<13>) );
	DFFPOSX1 DFFPOSX1_975 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4036), .Q(dp.rf.rf_8_<14>) );
	DFFPOSX1 DFFPOSX1_976 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4037), .Q(dp.rf.rf_8_<15>) );
	DFFPOSX1 DFFPOSX1_977 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4038), .Q(dp.rf.rf_8_<16>) );
	DFFPOSX1 DFFPOSX1_978 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4039), .Q(dp.rf.rf_8_<17>) );
	DFFPOSX1 DFFPOSX1_979 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4040), .Q(dp.rf.rf_8_<18>) );
	DFFPOSX1 DFFPOSX1_980 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4041), .Q(dp.rf.rf_8_<19>) );
	DFFPOSX1 DFFPOSX1_981 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4042), .Q(dp.rf.rf_8_<20>) );
	DFFPOSX1 DFFPOSX1_982 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4043), .Q(dp.rf.rf_8_<21>) );
	DFFPOSX1 DFFPOSX1_983 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4044), .Q(dp.rf.rf_8_<22>) );
	DFFPOSX1 DFFPOSX1_984 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4045), .Q(dp.rf.rf_8_<23>) );
	DFFPOSX1 DFFPOSX1_985 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4046), .Q(dp.rf.rf_8_<24>) );
	DFFPOSX1 DFFPOSX1_986 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4047), .Q(dp.rf.rf_8_<25>) );
	DFFPOSX1 DFFPOSX1_987 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4048), .Q(dp.rf.rf_8_<26>) );
	DFFPOSX1 DFFPOSX1_988 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4049), .Q(dp.rf.rf_8_<27>) );
	DFFPOSX1 DFFPOSX1_989 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4050), .Q(dp.rf.rf_8_<28>) );
	DFFPOSX1 DFFPOSX1_990 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4051), .Q(dp.rf.rf_8_<29>) );
	DFFPOSX1 DFFPOSX1_991 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4052), .Q(dp.rf.rf_8_<30>) );
	DFFPOSX1 DFFPOSX1_992 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4053), .Q(dp.rf.rf_8_<31>) );
	DFFPOSX1 DFFPOSX1_993 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4054), .Q(dp.rf.rf_9_<0>) );
	DFFPOSX1 DFFPOSX1_994 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4055), .Q(dp.rf.rf_9_<1>) );
	DFFPOSX1 DFFPOSX1_995 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4056), .Q(dp.rf.rf_9_<2>) );
	DFFPOSX1 DFFPOSX1_996 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4057), .Q(dp.rf.rf_9_<3>) );
	DFFPOSX1 DFFPOSX1_997 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4058), .Q(dp.rf.rf_9_<4>) );
	DFFPOSX1 DFFPOSX1_998 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4059), .Q(dp.rf.rf_9_<5>) );
	DFFPOSX1 DFFPOSX1_999 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4060), .Q(dp.rf.rf_9_<6>) );
	DFFPOSX1 DFFPOSX1_1000 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4061), .Q(dp.rf.rf_9_<7>) );
	DFFPOSX1 DFFPOSX1_1001 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4062), .Q(dp.rf.rf_9_<8>) );
	DFFPOSX1 DFFPOSX1_1002 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4063), .Q(dp.rf.rf_9_<9>) );
	DFFPOSX1 DFFPOSX1_1003 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4064), .Q(dp.rf.rf_9_<10>) );
	DFFPOSX1 DFFPOSX1_1004 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4065), .Q(dp.rf.rf_9_<11>) );
	DFFPOSX1 DFFPOSX1_1005 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4066), .Q(dp.rf.rf_9_<12>) );
	DFFPOSX1 DFFPOSX1_1006 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4067), .Q(dp.rf.rf_9_<13>) );
	DFFPOSX1 DFFPOSX1_1007 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4068), .Q(dp.rf.rf_9_<14>) );
	DFFPOSX1 DFFPOSX1_1008 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4069), .Q(dp.rf.rf_9_<15>) );
	DFFPOSX1 DFFPOSX1_1009 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4070), .Q(dp.rf.rf_9_<16>) );
	DFFPOSX1 DFFPOSX1_1010 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4071), .Q(dp.rf.rf_9_<17>) );
	DFFPOSX1 DFFPOSX1_1011 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4072), .Q(dp.rf.rf_9_<18>) );
	DFFPOSX1 DFFPOSX1_1012 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4073), .Q(dp.rf.rf_9_<19>) );
	DFFPOSX1 DFFPOSX1_1013 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4074), .Q(dp.rf.rf_9_<20>) );
	DFFPOSX1 DFFPOSX1_1014 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4075), .Q(dp.rf.rf_9_<21>) );
	DFFPOSX1 DFFPOSX1_1015 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4076), .Q(dp.rf.rf_9_<22>) );
	DFFPOSX1 DFFPOSX1_1016 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4077), .Q(dp.rf.rf_9_<23>) );
	DFFPOSX1 DFFPOSX1_1017 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4078), .Q(dp.rf.rf_9_<24>) );
	DFFPOSX1 DFFPOSX1_1018 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4079), .Q(dp.rf.rf_9_<25>) );
	DFFPOSX1 DFFPOSX1_1019 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4080), .Q(dp.rf.rf_9_<26>) );
	DFFPOSX1 DFFPOSX1_1020 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4081), .Q(dp.rf.rf_9_<27>) );
	DFFPOSX1 DFFPOSX1_1021 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4082), .Q(dp.rf.rf_9_<28>) );
	DFFPOSX1 DFFPOSX1_1022 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4083), .Q(dp.rf.rf_9_<29>) );
	DFFPOSX1 DFFPOSX1_1023 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4084), .Q(dp.rf.rf_9_<30>) );
	DFFPOSX1 DFFPOSX1_1024 ( .gnd(gnd), .vdd(vdd), .CLK(clk), .D(dp.rf._abc_6362_n4085), .Q(dp.rf.rf_9_<31>) );
	NAND2X1 NAND2X1_7841 ( .gnd(gnd), .vdd(vdd), .A(instr[0]), .B(alusrc), .Y(dp.srcbmux._abc_6353_n97) );
	INVX8 INVX8_47 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .Y(dp.srcbmux._abc_6353_n98) );
	NAND2X1 NAND2X1_7842 ( .gnd(gnd), .vdd(vdd), .A(writedata_0__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n99) );
	NAND2X1 NAND2X1_7843 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n97), .B(dp.srcbmux._abc_6353_n99), .Y(dp.srcb_0_) );
	NAND2X1 NAND2X1_7844 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[1]), .Y(dp.srcbmux._abc_6353_n101) );
	NAND2X1 NAND2X1_7845 ( .gnd(gnd), .vdd(vdd), .A(writedata_1__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n102) );
	NAND2X1 NAND2X1_7846 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n101), .B(dp.srcbmux._abc_6353_n102), .Y(dp.srcb_1_) );
	NAND2X1 NAND2X1_7847 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[2]), .Y(dp.srcbmux._abc_6353_n104) );
	NAND2X1 NAND2X1_7848 ( .gnd(gnd), .vdd(vdd), .A(writedata_2__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n105) );
	NAND2X1 NAND2X1_7849 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n104), .B(dp.srcbmux._abc_6353_n105), .Y(dp.srcb_2_) );
	NAND2X1 NAND2X1_7850 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[3]), .Y(dp.srcbmux._abc_6353_n107) );
	NAND2X1 NAND2X1_7851 ( .gnd(gnd), .vdd(vdd), .A(writedata_3__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n108) );
	NAND2X1 NAND2X1_7852 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n107), .B(dp.srcbmux._abc_6353_n108), .Y(dp.srcb_3_) );
	NAND2X1 NAND2X1_7853 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[4]), .Y(dp.srcbmux._abc_6353_n110) );
	NAND2X1 NAND2X1_7854 ( .gnd(gnd), .vdd(vdd), .A(writedata_4__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n111) );
	NAND2X1 NAND2X1_7855 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n110), .B(dp.srcbmux._abc_6353_n111), .Y(dp.srcb_4_) );
	NAND2X1 NAND2X1_7856 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[5]), .Y(dp.srcbmux._abc_6353_n113) );
	NAND2X1 NAND2X1_7857 ( .gnd(gnd), .vdd(vdd), .A(writedata_5__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n114) );
	NAND2X1 NAND2X1_7858 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n113), .B(dp.srcbmux._abc_6353_n114), .Y(dp.srcb_5_) );
	NAND2X1 NAND2X1_7859 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[6]), .Y(dp.srcbmux._abc_6353_n116) );
	NAND2X1 NAND2X1_7860 ( .gnd(gnd), .vdd(vdd), .A(writedata_6__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n117) );
	NAND2X1 NAND2X1_7861 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n116), .B(dp.srcbmux._abc_6353_n117), .Y(dp.srcb_6_) );
	NAND2X1 NAND2X1_7862 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[7]), .Y(dp.srcbmux._abc_6353_n119) );
	NAND2X1 NAND2X1_7863 ( .gnd(gnd), .vdd(vdd), .A(writedata_7__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n120) );
	NAND2X1 NAND2X1_7864 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n119), .B(dp.srcbmux._abc_6353_n120), .Y(dp.srcb_7_) );
	NAND2X1 NAND2X1_7865 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[8]), .Y(dp.srcbmux._abc_6353_n122) );
	NAND2X1 NAND2X1_7866 ( .gnd(gnd), .vdd(vdd), .A(writedata_8__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n123) );
	NAND2X1 NAND2X1_7867 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n122), .B(dp.srcbmux._abc_6353_n123), .Y(dp.srcb_8_) );
	NAND2X1 NAND2X1_7868 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[9]), .Y(dp.srcbmux._abc_6353_n125) );
	NAND2X1 NAND2X1_7869 ( .gnd(gnd), .vdd(vdd), .A(writedata_9__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n126) );
	NAND2X1 NAND2X1_7870 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n125), .B(dp.srcbmux._abc_6353_n126), .Y(dp.srcb_9_) );
	NAND2X1 NAND2X1_7871 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[10]), .Y(dp.srcbmux._abc_6353_n128) );
	NAND2X1 NAND2X1_7872 ( .gnd(gnd), .vdd(vdd), .A(writedata_10__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n129) );
	NAND2X1 NAND2X1_7873 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n128), .B(dp.srcbmux._abc_6353_n129), .Y(dp.srcb_10_) );
	NAND2X1 NAND2X1_7874 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[11]), .Y(dp.srcbmux._abc_6353_n131) );
	NAND2X1 NAND2X1_7875 ( .gnd(gnd), .vdd(vdd), .A(writedata_11__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n132) );
	NAND2X1 NAND2X1_7876 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n131), .B(dp.srcbmux._abc_6353_n132), .Y(dp.srcb_11_) );
	NAND2X1 NAND2X1_7877 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[12]), .Y(dp.srcbmux._abc_6353_n134) );
	NAND2X1 NAND2X1_7878 ( .gnd(gnd), .vdd(vdd), .A(writedata_12__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n135) );
	NAND2X1 NAND2X1_7879 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n134), .B(dp.srcbmux._abc_6353_n135), .Y(dp.srcb_12_) );
	NAND2X1 NAND2X1_7880 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[13]), .Y(dp.srcbmux._abc_6353_n137) );
	NAND2X1 NAND2X1_7881 ( .gnd(gnd), .vdd(vdd), .A(writedata_13__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n138) );
	NAND2X1 NAND2X1_7882 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n137), .B(dp.srcbmux._abc_6353_n138), .Y(dp.srcb_13_) );
	NAND2X1 NAND2X1_7883 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[14]), .Y(dp.srcbmux._abc_6353_n140) );
	NAND2X1 NAND2X1_7884 ( .gnd(gnd), .vdd(vdd), .A(writedata_14__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n141) );
	NAND2X1 NAND2X1_7885 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n140), .B(dp.srcbmux._abc_6353_n141), .Y(dp.srcb_14_) );
	NAND2X1 NAND2X1_7886 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n143) );
	NAND2X1 NAND2X1_7887 ( .gnd(gnd), .vdd(vdd), .A(writedata_15__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n144) );
	NAND2X1 NAND2X1_7888 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n143), .B(dp.srcbmux._abc_6353_n144), .Y(dp.srcb_15_) );
	NAND2X1 NAND2X1_7889 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n146) );
	NAND2X1 NAND2X1_7890 ( .gnd(gnd), .vdd(vdd), .A(writedata_16__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n147) );
	NAND2X1 NAND2X1_7891 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n146), .B(dp.srcbmux._abc_6353_n147), .Y(dp.srcb_16_) );
	NAND2X1 NAND2X1_7892 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n149) );
	NAND2X1 NAND2X1_7893 ( .gnd(gnd), .vdd(vdd), .A(writedata_17__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n150) );
	NAND2X1 NAND2X1_7894 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n149), .B(dp.srcbmux._abc_6353_n150), .Y(dp.srcb_17_) );
	NAND2X1 NAND2X1_7895 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n152) );
	NAND2X1 NAND2X1_7896 ( .gnd(gnd), .vdd(vdd), .A(writedata_18__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n153) );
	NAND2X1 NAND2X1_7897 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n152), .B(dp.srcbmux._abc_6353_n153), .Y(dp.srcb_18_) );
	NAND2X1 NAND2X1_7898 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n155) );
	NAND2X1 NAND2X1_7899 ( .gnd(gnd), .vdd(vdd), .A(writedata_19__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n156) );
	NAND2X1 NAND2X1_7900 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n155), .B(dp.srcbmux._abc_6353_n156), .Y(dp.srcb_19_) );
	NAND2X1 NAND2X1_7901 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n158) );
	NAND2X1 NAND2X1_7902 ( .gnd(gnd), .vdd(vdd), .A(writedata_20__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n159) );
	NAND2X1 NAND2X1_7903 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n158), .B(dp.srcbmux._abc_6353_n159), .Y(dp.srcb_20_) );
	NAND2X1 NAND2X1_7904 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n161) );
	NAND2X1 NAND2X1_7905 ( .gnd(gnd), .vdd(vdd), .A(writedata_21__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n162) );
	NAND2X1 NAND2X1_7906 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n161), .B(dp.srcbmux._abc_6353_n162), .Y(dp.srcb_21_) );
	NAND2X1 NAND2X1_7907 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n164) );
	NAND2X1 NAND2X1_7908 ( .gnd(gnd), .vdd(vdd), .A(writedata_22__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n165) );
	NAND2X1 NAND2X1_7909 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n164), .B(dp.srcbmux._abc_6353_n165), .Y(dp.srcb_22_) );
	NAND2X1 NAND2X1_7910 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n167) );
	NAND2X1 NAND2X1_7911 ( .gnd(gnd), .vdd(vdd), .A(writedata_23__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n168) );
	NAND2X1 NAND2X1_7912 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n167), .B(dp.srcbmux._abc_6353_n168), .Y(dp.srcb_23_) );
	NAND2X1 NAND2X1_7913 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n170) );
	NAND2X1 NAND2X1_7914 ( .gnd(gnd), .vdd(vdd), .A(writedata_24__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n171) );
	NAND2X1 NAND2X1_7915 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n170), .B(dp.srcbmux._abc_6353_n171), .Y(dp.srcb_24_) );
	NAND2X1 NAND2X1_7916 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n173) );
	NAND2X1 NAND2X1_7917 ( .gnd(gnd), .vdd(vdd), .A(writedata_25__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n174) );
	NAND2X1 NAND2X1_7918 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n173), .B(dp.srcbmux._abc_6353_n174), .Y(dp.srcb_25_) );
	NAND2X1 NAND2X1_7919 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n176) );
	NAND2X1 NAND2X1_7920 ( .gnd(gnd), .vdd(vdd), .A(writedata_26__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n177) );
	NAND2X1 NAND2X1_7921 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n176), .B(dp.srcbmux._abc_6353_n177), .Y(dp.srcb_26_) );
	NAND2X1 NAND2X1_7922 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n179) );
	NAND2X1 NAND2X1_7923 ( .gnd(gnd), .vdd(vdd), .A(writedata_27__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n180) );
	NAND2X1 NAND2X1_7924 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n179), .B(dp.srcbmux._abc_6353_n180), .Y(dp.srcb_27_) );
	NAND2X1 NAND2X1_7925 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n182) );
	NAND2X1 NAND2X1_7926 ( .gnd(gnd), .vdd(vdd), .A(writedata_28__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n183) );
	NAND2X1 NAND2X1_7927 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n182), .B(dp.srcbmux._abc_6353_n183), .Y(dp.srcb_28_) );
	NAND2X1 NAND2X1_7928 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n185) );
	NAND2X1 NAND2X1_7929 ( .gnd(gnd), .vdd(vdd), .A(writedata_29__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n186) );
	NAND2X1 NAND2X1_7930 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n185), .B(dp.srcbmux._abc_6353_n186), .Y(dp.srcb_29_) );
	NAND2X1 NAND2X1_7931 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n188) );
	NAND2X1 NAND2X1_7932 ( .gnd(gnd), .vdd(vdd), .A(writedata_30__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n189) );
	NAND2X1 NAND2X1_7933 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n188), .B(dp.srcbmux._abc_6353_n189), .Y(dp.srcb_30_) );
	NAND2X1 NAND2X1_7934 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .B(instr[15]), .Y(dp.srcbmux._abc_6353_n191) );
	NAND2X1 NAND2X1_7935 ( .gnd(gnd), .vdd(vdd), .A(writedata_31__RAW), .B(dp.srcbmux._abc_6353_n98), .Y(dp.srcbmux._abc_6353_n192) );
	NAND2X1 NAND2X1_7936 ( .gnd(gnd), .vdd(vdd), .A(dp.srcbmux._abc_6353_n191), .B(dp.srcbmux._abc_6353_n192), .Y(dp.srcb_31_) );
	NAND2X1 NAND2X1_7937 ( .gnd(gnd), .vdd(vdd), .A(instr[11]), .B(c.aluop_1_), .Y(dp.wrmux._abc_6354_n16) );
	INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_1_), .Y(dp.wrmux._abc_6354_n17) );
	NAND2X1 NAND2X1_7938 ( .gnd(gnd), .vdd(vdd), .A(instr[16]), .B(dp.wrmux._abc_6354_n17), .Y(dp.wrmux._abc_6354_n18) );
	NAND2X1 NAND2X1_7939 ( .gnd(gnd), .vdd(vdd), .A(dp.wrmux._abc_6354_n16), .B(dp.wrmux._abc_6354_n18), .Y(dp.writereg_0_) );
	NAND2X1 NAND2X1_7940 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_1_), .B(instr[12]), .Y(dp.wrmux._abc_6354_n20) );
	NAND2X1 NAND2X1_7941 ( .gnd(gnd), .vdd(vdd), .A(instr[17]), .B(dp.wrmux._abc_6354_n17), .Y(dp.wrmux._abc_6354_n21) );
	NAND2X1 NAND2X1_7942 ( .gnd(gnd), .vdd(vdd), .A(dp.wrmux._abc_6354_n20), .B(dp.wrmux._abc_6354_n21), .Y(dp.writereg_1_) );
	NAND2X1 NAND2X1_7943 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_1_), .B(instr[13]), .Y(dp.wrmux._abc_6354_n23) );
	NAND2X1 NAND2X1_7944 ( .gnd(gnd), .vdd(vdd), .A(instr[18]), .B(dp.wrmux._abc_6354_n17), .Y(dp.wrmux._abc_6354_n24) );
	NAND2X1 NAND2X1_7945 ( .gnd(gnd), .vdd(vdd), .A(dp.wrmux._abc_6354_n23), .B(dp.wrmux._abc_6354_n24), .Y(dp.writereg_2_) );
	NAND2X1 NAND2X1_7946 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_1_), .B(instr[14]), .Y(dp.wrmux._abc_6354_n26) );
	NAND2X1 NAND2X1_7947 ( .gnd(gnd), .vdd(vdd), .A(instr[19]), .B(dp.wrmux._abc_6354_n17), .Y(dp.wrmux._abc_6354_n27) );
	NAND2X1 NAND2X1_7948 ( .gnd(gnd), .vdd(vdd), .A(dp.wrmux._abc_6354_n26), .B(dp.wrmux._abc_6354_n27), .Y(dp.writereg_3_) );
	NAND2X1 NAND2X1_7949 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_1_), .B(instr[15]), .Y(dp.wrmux._abc_6354_n29) );
	NAND2X1 NAND2X1_7950 ( .gnd(gnd), .vdd(vdd), .A(instr[20]), .B(dp.wrmux._abc_6354_n17), .Y(dp.wrmux._abc_6354_n30) );
	NAND2X1 NAND2X1_7951 ( .gnd(gnd), .vdd(vdd), .A(dp.wrmux._abc_6354_n29), .B(dp.wrmux._abc_6354_n30), .Y(dp.writereg_4_) );
	BUFX2 BUFX2_98 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_0_), .Y(c.branch) );
	BUFX2 BUFX2_99 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_0_), .Y(c.md.controls_0_) );
	BUFX2 BUFX2_100 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_1_), .Y(c.md.controls_1_) );
	BUFX2 BUFX2_101 ( .gnd(gnd), .vdd(vdd), .A(memwrite_RAW), .Y(c.md.controls_4_) );
	BUFX2 BUFX2_102 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_0_), .Y(c.md.controls_5_) );
	BUFX2 BUFX2_103 ( .gnd(gnd), .vdd(vdd), .A(alusrc), .Y(c.md.controls_6_) );
	BUFX2 BUFX2_104 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_1_), .Y(c.md.controls_7_) );
	BUFX2 BUFX2_105 ( .gnd(gnd), .vdd(vdd), .A(instr[0]), .Y(dp.signimm_0_) );
	BUFX2 BUFX2_106 ( .gnd(gnd), .vdd(vdd), .A(instr[1]), .Y(dp.signimm_1_) );
	BUFX2 BUFX2_107 ( .gnd(gnd), .vdd(vdd), .A(instr[2]), .Y(dp.signimm_2_) );
	BUFX2 BUFX2_108 ( .gnd(gnd), .vdd(vdd), .A(instr[3]), .Y(dp.signimm_3_) );
	BUFX2 BUFX2_109 ( .gnd(gnd), .vdd(vdd), .A(instr[4]), .Y(dp.signimm_4_) );
	BUFX2 BUFX2_110 ( .gnd(gnd), .vdd(vdd), .A(instr[5]), .Y(dp.signimm_5_) );
	BUFX2 BUFX2_111 ( .gnd(gnd), .vdd(vdd), .A(instr[6]), .Y(dp.signimm_6_) );
	BUFX2 BUFX2_112 ( .gnd(gnd), .vdd(vdd), .A(instr[7]), .Y(dp.signimm_7_) );
	BUFX2 BUFX2_113 ( .gnd(gnd), .vdd(vdd), .A(instr[8]), .Y(dp.signimm_8_) );
	BUFX2 BUFX2_114 ( .gnd(gnd), .vdd(vdd), .A(instr[9]), .Y(dp.signimm_9_) );
	BUFX2 BUFX2_115 ( .gnd(gnd), .vdd(vdd), .A(instr[10]), .Y(dp.signimm_10_) );
	BUFX2 BUFX2_116 ( .gnd(gnd), .vdd(vdd), .A(instr[11]), .Y(dp.signimm_11_) );
	BUFX2 BUFX2_117 ( .gnd(gnd), .vdd(vdd), .A(instr[12]), .Y(dp.signimm_12_) );
	BUFX2 BUFX2_118 ( .gnd(gnd), .vdd(vdd), .A(instr[13]), .Y(dp.signimm_13_) );
	BUFX2 BUFX2_119 ( .gnd(gnd), .vdd(vdd), .A(instr[14]), .Y(dp.signimm_14_) );
	BUFX2 BUFX2_120 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_15_) );
	BUFX2 BUFX2_121 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_16_) );
	BUFX2 BUFX2_122 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_17_) );
	BUFX2 BUFX2_123 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_18_) );
	BUFX2 BUFX2_124 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_19_) );
	BUFX2 BUFX2_125 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_20_) );
	BUFX2 BUFX2_126 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_21_) );
	BUFX2 BUFX2_127 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_22_) );
	BUFX2 BUFX2_128 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_23_) );
	BUFX2 BUFX2_129 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_24_) );
	BUFX2 BUFX2_130 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_25_) );
	BUFX2 BUFX2_131 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_26_) );
	BUFX2 BUFX2_132 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_27_) );
	BUFX2 BUFX2_133 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_28_) );
	BUFX2 BUFX2_134 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_29_) );
	BUFX2 BUFX2_135 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_30_) );
	BUFX2 BUFX2_136 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimm_31_) );
	BUFX2 BUFX2_137 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(dp.signimmsh_0_) );
	BUFX2 BUFX2_138 ( .gnd(gnd), .vdd(vdd), .A(gnd), .Y(dp.signimmsh_1_) );
	BUFX2 BUFX2_139 ( .gnd(gnd), .vdd(vdd), .A(instr[0]), .Y(dp.signimmsh_2_) );
	BUFX2 BUFX2_140 ( .gnd(gnd), .vdd(vdd), .A(instr[1]), .Y(dp.signimmsh_3_) );
	BUFX2 BUFX2_141 ( .gnd(gnd), .vdd(vdd), .A(instr[2]), .Y(dp.signimmsh_4_) );
	BUFX2 BUFX2_142 ( .gnd(gnd), .vdd(vdd), .A(instr[3]), .Y(dp.signimmsh_5_) );
	BUFX2 BUFX2_143 ( .gnd(gnd), .vdd(vdd), .A(instr[4]), .Y(dp.signimmsh_6_) );
	BUFX2 BUFX2_144 ( .gnd(gnd), .vdd(vdd), .A(instr[5]), .Y(dp.signimmsh_7_) );
	BUFX2 BUFX2_145 ( .gnd(gnd), .vdd(vdd), .A(instr[6]), .Y(dp.signimmsh_8_) );
	BUFX2 BUFX2_146 ( .gnd(gnd), .vdd(vdd), .A(instr[7]), .Y(dp.signimmsh_9_) );
	BUFX2 BUFX2_147 ( .gnd(gnd), .vdd(vdd), .A(instr[8]), .Y(dp.signimmsh_10_) );
	BUFX2 BUFX2_148 ( .gnd(gnd), .vdd(vdd), .A(instr[9]), .Y(dp.signimmsh_11_) );
	BUFX2 BUFX2_149 ( .gnd(gnd), .vdd(vdd), .A(instr[10]), .Y(dp.signimmsh_12_) );
	BUFX2 BUFX2_150 ( .gnd(gnd), .vdd(vdd), .A(instr[11]), .Y(dp.signimmsh_13_) );
	BUFX2 BUFX2_151 ( .gnd(gnd), .vdd(vdd), .A(instr[12]), .Y(dp.signimmsh_14_) );
	BUFX2 BUFX2_152 ( .gnd(gnd), .vdd(vdd), .A(instr[13]), .Y(dp.signimmsh_15_) );
	BUFX2 BUFX2_153 ( .gnd(gnd), .vdd(vdd), .A(instr[14]), .Y(dp.signimmsh_16_) );
	BUFX2 BUFX2_154 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_17_) );
	BUFX2 BUFX2_155 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_18_) );
	BUFX2 BUFX2_156 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_19_) );
	BUFX2 BUFX2_157 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_20_) );
	BUFX2 BUFX2_158 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_21_) );
	BUFX2 BUFX2_159 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_22_) );
	BUFX2 BUFX2_160 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_23_) );
	BUFX2 BUFX2_161 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_24_) );
	BUFX2 BUFX2_162 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_25_) );
	BUFX2 BUFX2_163 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_26_) );
	BUFX2 BUFX2_164 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_27_) );
	BUFX2 BUFX2_165 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_28_) );
	BUFX2 BUFX2_166 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_29_) );
	BUFX2 BUFX2_167 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_30_) );
	BUFX2 BUFX2_168 ( .gnd(gnd), .vdd(vdd), .A(instr[15]), .Y(dp.signimmsh_31_) );
	BUFX2 BUFX2_169 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_2_), .Y(jump) );
	BUFX2 BUFX2_170 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_3_), .Y(memtoreg) );
	BUFX2 BUFX2_171 ( .gnd(gnd), .vdd(vdd), .A(c.aluop_1_), .Y(regdst) );
	BUFX2 BUFX2_172 ( .gnd(gnd), .vdd(vdd), .A(c.md.controls_8_), .Y(regwrite) );
endmodule
